// -----------------------------------------------------------------------------
// Title   : Pipeline ROM 1A (Pipeline/roms/Pipe1A.v)
// Create  : Thu, Dec 22, 2022  5:55:34 PM
//
// Name    : JAM-1 8-bit Pipelined CPU in Verilog
// Author  : George Smart, M1GEO.  https://www.george-smart.co.uk
// GitHub  : https://github.com/m1geo/JamesSharmanPipelinedCPU
// CPU Dsn : James Sharman; Video Series => https://youtu.be/3iHag4k4yEg
//
// Desc.   : Pipeline ROM 1A
// -----------------------------------------------------------------------------

module pipeline_rom_1a
(
    input         clk,
    input         en, // active high
    input  [14:0] addr,
    output  [7:0] dout
);

    (*rom_style = "block" *) reg [7:0] d;

    always @ (posedge clk) begin
        if (en)
            case(addr)
                15'h0000: d <= 8'hC0; 15'h0001: d <= 8'hC0; 15'h0002: d <= 8'hC0; 15'h0003: d <= 8'hC0;
                15'h0004: d <= 8'hC0; 15'h0005: d <= 8'hC0; 15'h0006: d <= 8'hC0; 15'h0007: d <= 8'hC0;
                15'h0008: d <= 8'hC0; 15'h0009: d <= 8'hC0; 15'h000A: d <= 8'hC0; 15'h000B: d <= 8'hC0;
                15'h000C: d <= 8'hC0; 15'h000D: d <= 8'hC0; 15'h000E: d <= 8'hC0; 15'h000F: d <= 8'hC0;
                15'h0010: d <= 8'hC0; 15'h0011: d <= 8'hC0; 15'h0012: d <= 8'hC0; 15'h0013: d <= 8'hC0;
                15'h0014: d <= 8'hC0; 15'h0015: d <= 8'hC0; 15'h0016: d <= 8'hC0; 15'h0017: d <= 8'hC0;
                15'h0018: d <= 8'hC0; 15'h0019: d <= 8'hC0; 15'h001A: d <= 8'hC0; 15'h001B: d <= 8'hC0;
                15'h001C: d <= 8'hC0; 15'h001D: d <= 8'hC0; 15'h001E: d <= 8'hC0; 15'h001F: d <= 8'hC0;
                15'h0020: d <= 8'hC0; 15'h0021: d <= 8'hC0; 15'h0022: d <= 8'hC0; 15'h0023: d <= 8'hC0;
                15'h0024: d <= 8'hC0; 15'h0025: d <= 8'hC0; 15'h0026: d <= 8'hC0; 15'h0027: d <= 8'hC0;
                15'h0028: d <= 8'hC0; 15'h0029: d <= 8'hC0; 15'h002A: d <= 8'hC0; 15'h002B: d <= 8'hC0;
                15'h002C: d <= 8'hC0; 15'h002D: d <= 8'hC0; 15'h002E: d <= 8'hC0; 15'h002F: d <= 8'hC0;
                15'h0030: d <= 8'hC0; 15'h0031: d <= 8'hC0; 15'h0032: d <= 8'hC0; 15'h0033: d <= 8'hC0;
                15'h0034: d <= 8'hC0; 15'h0035: d <= 8'hC0; 15'h0036: d <= 8'hC0; 15'h0037: d <= 8'hC0;
                15'h0038: d <= 8'hC0; 15'h0039: d <= 8'hC0; 15'h003A: d <= 8'hC0; 15'h003B: d <= 8'hC0;
                15'h003C: d <= 8'hC0; 15'h003D: d <= 8'hC0; 15'h003E: d <= 8'hC0; 15'h003F: d <= 8'hC0;
                15'h0040: d <= 8'hC0; 15'h0041: d <= 8'hC0; 15'h0042: d <= 8'hC0; 15'h0043: d <= 8'hC0;
                15'h0044: d <= 8'hC0; 15'h0045: d <= 8'hC0; 15'h0046: d <= 8'hC0; 15'h0047: d <= 8'hC0;
                15'h0048: d <= 8'hC0; 15'h0049: d <= 8'hC0; 15'h004A: d <= 8'hC0; 15'h004B: d <= 8'hC0;
                15'h004C: d <= 8'hC0; 15'h004D: d <= 8'hC0; 15'h004E: d <= 8'hC0; 15'h004F: d <= 8'hC0;
                15'h0050: d <= 8'hC0; 15'h0051: d <= 8'hC0; 15'h0052: d <= 8'hC0; 15'h0053: d <= 8'hC0;
                15'h0054: d <= 8'hC0; 15'h0055: d <= 8'hC0; 15'h0056: d <= 8'hC0; 15'h0057: d <= 8'hC0;
                15'h0058: d <= 8'hC0; 15'h0059: d <= 8'hC0; 15'h005A: d <= 8'hC0; 15'h005B: d <= 8'hC0;
                15'h005C: d <= 8'hC0; 15'h005D: d <= 8'hC0; 15'h005E: d <= 8'hC0; 15'h005F: d <= 8'hC0;
                15'h0060: d <= 8'hC0; 15'h0061: d <= 8'hC0; 15'h0062: d <= 8'hC0; 15'h0063: d <= 8'hC0;
                15'h0064: d <= 8'hC0; 15'h0065: d <= 8'hC0; 15'h0066: d <= 8'hC0; 15'h0067: d <= 8'hC0;
                15'h0068: d <= 8'hC0; 15'h0069: d <= 8'hC0; 15'h006A: d <= 8'hC0; 15'h006B: d <= 8'hC0;
                15'h006C: d <= 8'hC0; 15'h006D: d <= 8'hC0; 15'h006E: d <= 8'hC0; 15'h006F: d <= 8'hC0;
                15'h0070: d <= 8'hC0; 15'h0071: d <= 8'hC0; 15'h0072: d <= 8'hC0; 15'h0073: d <= 8'hC0;
                15'h0074: d <= 8'hC0; 15'h0075: d <= 8'hC0; 15'h0076: d <= 8'hC0; 15'h0077: d <= 8'hC0;
                15'h0078: d <= 8'hC0; 15'h0079: d <= 8'hC0; 15'h007A: d <= 8'hC0; 15'h007B: d <= 8'hC0;
                15'h007C: d <= 8'hC0; 15'h007D: d <= 8'hC0; 15'h007E: d <= 8'hC0; 15'h007F: d <= 8'hC0;
                15'h0080: d <= 8'hC0; 15'h0081: d <= 8'hC0; 15'h0082: d <= 8'hC0; 15'h0083: d <= 8'hC0;
                15'h0084: d <= 8'hC0; 15'h0085: d <= 8'hC0; 15'h0086: d <= 8'hC0; 15'h0087: d <= 8'hC0;
                15'h0088: d <= 8'hC0; 15'h0089: d <= 8'hC0; 15'h008A: d <= 8'hC0; 15'h008B: d <= 8'hC0;
                15'h008C: d <= 8'hC0; 15'h008D: d <= 8'hC0; 15'h008E: d <= 8'hC0; 15'h008F: d <= 8'hC0;
                15'h0090: d <= 8'hC0; 15'h0091: d <= 8'hC0; 15'h0092: d <= 8'hC0; 15'h0093: d <= 8'hC0;
                15'h0094: d <= 8'hC0; 15'h0095: d <= 8'hC0; 15'h0096: d <= 8'hC0; 15'h0097: d <= 8'hC0;
                15'h0098: d <= 8'hC0; 15'h0099: d <= 8'hC0; 15'h009A: d <= 8'hC0; 15'h009B: d <= 8'hC0;
                15'h009C: d <= 8'hC0; 15'h009D: d <= 8'hC0; 15'h009E: d <= 8'hC0; 15'h009F: d <= 8'hC0;
                15'h00A0: d <= 8'hC0; 15'h00A1: d <= 8'hC0; 15'h00A2: d <= 8'hC0; 15'h00A3: d <= 8'hC0;
                15'h00A4: d <= 8'hC0; 15'h00A5: d <= 8'hC0; 15'h00A6: d <= 8'hC0; 15'h00A7: d <= 8'hC0;
                15'h00A8: d <= 8'hC0; 15'h00A9: d <= 8'hC0; 15'h00AA: d <= 8'hC0; 15'h00AB: d <= 8'hC0;
                15'h00AC: d <= 8'hC0; 15'h00AD: d <= 8'hC0; 15'h00AE: d <= 8'hC0; 15'h00AF: d <= 8'hC0;
                15'h00B0: d <= 8'hC0; 15'h00B1: d <= 8'hC0; 15'h00B2: d <= 8'hC0; 15'h00B3: d <= 8'hC0;
                15'h00B4: d <= 8'hC0; 15'h00B5: d <= 8'hC0; 15'h00B6: d <= 8'hC0; 15'h00B7: d <= 8'hC0;
                15'h00B8: d <= 8'hC0; 15'h00B9: d <= 8'hC0; 15'h00BA: d <= 8'hC0; 15'h00BB: d <= 8'hC0;
                15'h00BC: d <= 8'hC0; 15'h00BD: d <= 8'hC0; 15'h00BE: d <= 8'hC0; 15'h00BF: d <= 8'hC0;
                15'h00C0: d <= 8'hC0; 15'h00C1: d <= 8'hC0; 15'h00C2: d <= 8'hC0; 15'h00C3: d <= 8'hC0;
                15'h00C4: d <= 8'hC0; 15'h00C5: d <= 8'hC0; 15'h00C6: d <= 8'hC0; 15'h00C7: d <= 8'hC0;
                15'h00C8: d <= 8'hC0; 15'h00C9: d <= 8'hC0; 15'h00CA: d <= 8'hC0; 15'h00CB: d <= 8'hC0;
                15'h00CC: d <= 8'hC0; 15'h00CD: d <= 8'hC0; 15'h00CE: d <= 8'hC0; 15'h00CF: d <= 8'hC0;
                15'h00D0: d <= 8'hC0; 15'h00D1: d <= 8'hC0; 15'h00D2: d <= 8'hC0; 15'h00D3: d <= 8'hC0;
                15'h00D4: d <= 8'hC0; 15'h00D5: d <= 8'hC0; 15'h00D6: d <= 8'hC0; 15'h00D7: d <= 8'hC0;
                15'h00D8: d <= 8'hC0; 15'h00D9: d <= 8'hC0; 15'h00DA: d <= 8'hC0; 15'h00DB: d <= 8'hC0;
                15'h00DC: d <= 8'hC0; 15'h00DD: d <= 8'hC0; 15'h00DE: d <= 8'hC0; 15'h00DF: d <= 8'hC0;
                15'h00E0: d <= 8'hC0; 15'h00E1: d <= 8'hC0; 15'h00E2: d <= 8'hC0; 15'h00E3: d <= 8'hC0;
                15'h00E4: d <= 8'hC0; 15'h00E5: d <= 8'hC0; 15'h00E6: d <= 8'hC0; 15'h00E7: d <= 8'hC0;
                15'h00E8: d <= 8'hC0; 15'h00E9: d <= 8'hC0; 15'h00EA: d <= 8'hC0; 15'h00EB: d <= 8'hC0;
                15'h00EC: d <= 8'hC0; 15'h00ED: d <= 8'hC0; 15'h00EE: d <= 8'hC0; 15'h00EF: d <= 8'hC0;
                15'h00F0: d <= 8'hC0; 15'h00F1: d <= 8'hC0; 15'h00F2: d <= 8'hC0; 15'h00F3: d <= 8'hC0;
                15'h00F4: d <= 8'hC0; 15'h00F5: d <= 8'hC0; 15'h00F6: d <= 8'hC0; 15'h00F7: d <= 8'hC0;
                15'h00F8: d <= 8'hC0; 15'h00F9: d <= 8'hC0; 15'h00FA: d <= 8'hC0; 15'h00FB: d <= 8'hC0;
                15'h00FC: d <= 8'hC0; 15'h00FD: d <= 8'hC0; 15'h00FE: d <= 8'hC0; 15'h00FF: d <= 8'hC0;
                15'h0100: d <= 8'hC0; 15'h0101: d <= 8'hC0; 15'h0102: d <= 8'hC0; 15'h0103: d <= 8'hC0;
                15'h0104: d <= 8'hC0; 15'h0105: d <= 8'hC0; 15'h0106: d <= 8'hC0; 15'h0107: d <= 8'hC0;
                15'h0108: d <= 8'hC0; 15'h0109: d <= 8'hC0; 15'h010A: d <= 8'hC0; 15'h010B: d <= 8'hC0;
                15'h010C: d <= 8'hC0; 15'h010D: d <= 8'hC0; 15'h010E: d <= 8'hC0; 15'h010F: d <= 8'hC0;
                15'h0110: d <= 8'hC0; 15'h0111: d <= 8'hC0; 15'h0112: d <= 8'hC0; 15'h0113: d <= 8'hC0;
                15'h0114: d <= 8'hC0; 15'h0115: d <= 8'hC0; 15'h0116: d <= 8'hC0; 15'h0117: d <= 8'hC0;
                15'h0118: d <= 8'hC0; 15'h0119: d <= 8'hC0; 15'h011A: d <= 8'hC0; 15'h011B: d <= 8'hC0;
                15'h011C: d <= 8'hC0; 15'h011D: d <= 8'hC0; 15'h011E: d <= 8'hC0; 15'h011F: d <= 8'hC0;
                15'h0120: d <= 8'hC0; 15'h0121: d <= 8'hC0; 15'h0122: d <= 8'hC0; 15'h0123: d <= 8'hC0;
                15'h0124: d <= 8'hC0; 15'h0125: d <= 8'hC0; 15'h0126: d <= 8'hC0; 15'h0127: d <= 8'hC0;
                15'h0128: d <= 8'hC0; 15'h0129: d <= 8'hC0; 15'h012A: d <= 8'hC0; 15'h012B: d <= 8'hC0;
                15'h012C: d <= 8'hC0; 15'h012D: d <= 8'hC0; 15'h012E: d <= 8'hC0; 15'h012F: d <= 8'hC0;
                15'h0130: d <= 8'hC0; 15'h0131: d <= 8'hC0; 15'h0132: d <= 8'hC0; 15'h0133: d <= 8'hC0;
                15'h0134: d <= 8'hC0; 15'h0135: d <= 8'hC0; 15'h0136: d <= 8'hC0; 15'h0137: d <= 8'hC0;
                15'h0138: d <= 8'hC0; 15'h0139: d <= 8'hC0; 15'h013A: d <= 8'hC0; 15'h013B: d <= 8'hC0;
                15'h013C: d <= 8'hC0; 15'h013D: d <= 8'hC0; 15'h013E: d <= 8'hC0; 15'h013F: d <= 8'hC0;
                15'h0140: d <= 8'hC0; 15'h0141: d <= 8'hC0; 15'h0142: d <= 8'hC0; 15'h0143: d <= 8'hC0;
                15'h0144: d <= 8'hC0; 15'h0145: d <= 8'hC0; 15'h0146: d <= 8'hC0; 15'h0147: d <= 8'hC0;
                15'h0148: d <= 8'hC0; 15'h0149: d <= 8'hC0; 15'h014A: d <= 8'hC0; 15'h014B: d <= 8'hC0;
                15'h014C: d <= 8'hC0; 15'h014D: d <= 8'hC0; 15'h014E: d <= 8'hC0; 15'h014F: d <= 8'hC0;
                15'h0150: d <= 8'hC0; 15'h0151: d <= 8'hC0; 15'h0152: d <= 8'hC0; 15'h0153: d <= 8'hC0;
                15'h0154: d <= 8'hC0; 15'h0155: d <= 8'hC0; 15'h0156: d <= 8'hC0; 15'h0157: d <= 8'hC0;
                15'h0158: d <= 8'hC0; 15'h0159: d <= 8'hC0; 15'h015A: d <= 8'hC0; 15'h015B: d <= 8'hC0;
                15'h015C: d <= 8'hC0; 15'h015D: d <= 8'hC0; 15'h015E: d <= 8'hC0; 15'h015F: d <= 8'hC0;
                15'h0160: d <= 8'hC0; 15'h0161: d <= 8'hC0; 15'h0162: d <= 8'hC0; 15'h0163: d <= 8'hC0;
                15'h0164: d <= 8'hC0; 15'h0165: d <= 8'hC0; 15'h0166: d <= 8'hC0; 15'h0167: d <= 8'hC0;
                15'h0168: d <= 8'hC0; 15'h0169: d <= 8'hC0; 15'h016A: d <= 8'hC0; 15'h016B: d <= 8'hC0;
                15'h016C: d <= 8'hC0; 15'h016D: d <= 8'hC0; 15'h016E: d <= 8'hC0; 15'h016F: d <= 8'hC0;
                15'h0170: d <= 8'hC0; 15'h0171: d <= 8'hC0; 15'h0172: d <= 8'hC0; 15'h0173: d <= 8'hC0;
                15'h0174: d <= 8'hC0; 15'h0175: d <= 8'hC0; 15'h0176: d <= 8'hC0; 15'h0177: d <= 8'hC0;
                15'h0178: d <= 8'hC0; 15'h0179: d <= 8'hC0; 15'h017A: d <= 8'hC0; 15'h017B: d <= 8'hC0;
                15'h017C: d <= 8'hC0; 15'h017D: d <= 8'hC0; 15'h017E: d <= 8'hC0; 15'h017F: d <= 8'hC0;
                15'h0180: d <= 8'hC0; 15'h0181: d <= 8'hC0; 15'h0182: d <= 8'hC0; 15'h0183: d <= 8'hC0;
                15'h0184: d <= 8'hC0; 15'h0185: d <= 8'hC0; 15'h0186: d <= 8'hC0; 15'h0187: d <= 8'hC0;
                15'h0188: d <= 8'hC0; 15'h0189: d <= 8'hC0; 15'h018A: d <= 8'hC0; 15'h018B: d <= 8'hC0;
                15'h018C: d <= 8'hC0; 15'h018D: d <= 8'hC0; 15'h018E: d <= 8'hC0; 15'h018F: d <= 8'hC0;
                15'h0190: d <= 8'hC0; 15'h0191: d <= 8'hC0; 15'h0192: d <= 8'hC0; 15'h0193: d <= 8'hC0;
                15'h0194: d <= 8'hC0; 15'h0195: d <= 8'hC0; 15'h0196: d <= 8'hC0; 15'h0197: d <= 8'hC0;
                15'h0198: d <= 8'hC0; 15'h0199: d <= 8'hC0; 15'h019A: d <= 8'hC0; 15'h019B: d <= 8'hC0;
                15'h019C: d <= 8'hC0; 15'h019D: d <= 8'hC0; 15'h019E: d <= 8'hC0; 15'h019F: d <= 8'hC0;
                15'h01A0: d <= 8'hC0; 15'h01A1: d <= 8'hC0; 15'h01A2: d <= 8'hC0; 15'h01A3: d <= 8'hC0;
                15'h01A4: d <= 8'hC0; 15'h01A5: d <= 8'hC0; 15'h01A6: d <= 8'hC0; 15'h01A7: d <= 8'hC0;
                15'h01A8: d <= 8'hC0; 15'h01A9: d <= 8'hC0; 15'h01AA: d <= 8'hC0; 15'h01AB: d <= 8'hC0;
                15'h01AC: d <= 8'hC0; 15'h01AD: d <= 8'hC0; 15'h01AE: d <= 8'hC0; 15'h01AF: d <= 8'hC0;
                15'h01B0: d <= 8'hC0; 15'h01B1: d <= 8'hC0; 15'h01B2: d <= 8'hC0; 15'h01B3: d <= 8'hC0;
                15'h01B4: d <= 8'hC0; 15'h01B5: d <= 8'hC0; 15'h01B6: d <= 8'hC0; 15'h01B7: d <= 8'hC0;
                15'h01B8: d <= 8'hC0; 15'h01B9: d <= 8'hC0; 15'h01BA: d <= 8'hC0; 15'h01BB: d <= 8'hC0;
                15'h01BC: d <= 8'hC0; 15'h01BD: d <= 8'hC0; 15'h01BE: d <= 8'hC0; 15'h01BF: d <= 8'hC0;
                15'h01C0: d <= 8'hC0; 15'h01C1: d <= 8'hC0; 15'h01C2: d <= 8'hC0; 15'h01C3: d <= 8'hC0;
                15'h01C4: d <= 8'hC0; 15'h01C5: d <= 8'hC0; 15'h01C6: d <= 8'hC0; 15'h01C7: d <= 8'hC0;
                15'h01C8: d <= 8'hC0; 15'h01C9: d <= 8'hC0; 15'h01CA: d <= 8'hC0; 15'h01CB: d <= 8'hC0;
                15'h01CC: d <= 8'hC0; 15'h01CD: d <= 8'hC0; 15'h01CE: d <= 8'hC0; 15'h01CF: d <= 8'hC0;
                15'h01D0: d <= 8'hC0; 15'h01D1: d <= 8'hC0; 15'h01D2: d <= 8'hC0; 15'h01D3: d <= 8'hC0;
                15'h01D4: d <= 8'hC0; 15'h01D5: d <= 8'hC0; 15'h01D6: d <= 8'hC0; 15'h01D7: d <= 8'hC0;
                15'h01D8: d <= 8'hC0; 15'h01D9: d <= 8'hC0; 15'h01DA: d <= 8'hC0; 15'h01DB: d <= 8'hC0;
                15'h01DC: d <= 8'hC0; 15'h01DD: d <= 8'hC0; 15'h01DE: d <= 8'hC0; 15'h01DF: d <= 8'hC0;
                15'h01E0: d <= 8'hC0; 15'h01E1: d <= 8'hC0; 15'h01E2: d <= 8'hC0; 15'h01E3: d <= 8'hC0;
                15'h01E4: d <= 8'hC0; 15'h01E5: d <= 8'hC0; 15'h01E6: d <= 8'hC0; 15'h01E7: d <= 8'hC0;
                15'h01E8: d <= 8'hC0; 15'h01E9: d <= 8'hC0; 15'h01EA: d <= 8'hC0; 15'h01EB: d <= 8'hC0;
                15'h01EC: d <= 8'hC0; 15'h01ED: d <= 8'hC0; 15'h01EE: d <= 8'hC0; 15'h01EF: d <= 8'hC0;
                15'h01F0: d <= 8'hC0; 15'h01F1: d <= 8'hC0; 15'h01F2: d <= 8'hC0; 15'h01F3: d <= 8'hC0;
                15'h01F4: d <= 8'hC0; 15'h01F5: d <= 8'hC0; 15'h01F6: d <= 8'hC0; 15'h01F7: d <= 8'hC0;
                15'h01F8: d <= 8'hC0; 15'h01F9: d <= 8'hC0; 15'h01FA: d <= 8'hC0; 15'h01FB: d <= 8'hC0;
                15'h01FC: d <= 8'hC0; 15'h01FD: d <= 8'hC0; 15'h01FE: d <= 8'hC0; 15'h01FF: d <= 8'hC0;
                15'h0200: d <= 8'hC0; 15'h0201: d <= 8'hC0; 15'h0202: d <= 8'hC0; 15'h0203: d <= 8'hC0;
                15'h0204: d <= 8'hC0; 15'h0205: d <= 8'hC0; 15'h0206: d <= 8'hC0; 15'h0207: d <= 8'hC0;
                15'h0208: d <= 8'hC0; 15'h0209: d <= 8'hC0; 15'h020A: d <= 8'hC0; 15'h020B: d <= 8'hC0;
                15'h020C: d <= 8'hC0; 15'h020D: d <= 8'hC0; 15'h020E: d <= 8'hC0; 15'h020F: d <= 8'hC0;
                15'h0210: d <= 8'hC0; 15'h0211: d <= 8'hC0; 15'h0212: d <= 8'hC0; 15'h0213: d <= 8'hC0;
                15'h0214: d <= 8'hC0; 15'h0215: d <= 8'hC0; 15'h0216: d <= 8'hC0; 15'h0217: d <= 8'hC0;
                15'h0218: d <= 8'hC0; 15'h0219: d <= 8'hC0; 15'h021A: d <= 8'hC0; 15'h021B: d <= 8'hC0;
                15'h021C: d <= 8'hC0; 15'h021D: d <= 8'hC0; 15'h021E: d <= 8'hC0; 15'h021F: d <= 8'hC0;
                15'h0220: d <= 8'hC0; 15'h0221: d <= 8'hC0; 15'h0222: d <= 8'hC0; 15'h0223: d <= 8'hC0;
                15'h0224: d <= 8'hC0; 15'h0225: d <= 8'hC0; 15'h0226: d <= 8'hC0; 15'h0227: d <= 8'hC0;
                15'h0228: d <= 8'hC0; 15'h0229: d <= 8'hC0; 15'h022A: d <= 8'hC0; 15'h022B: d <= 8'hC0;
                15'h022C: d <= 8'hC0; 15'h022D: d <= 8'hC0; 15'h022E: d <= 8'hC0; 15'h022F: d <= 8'hC0;
                15'h0230: d <= 8'hC0; 15'h0231: d <= 8'hC0; 15'h0232: d <= 8'hC0; 15'h0233: d <= 8'hC0;
                15'h0234: d <= 8'hC0; 15'h0235: d <= 8'hC0; 15'h0236: d <= 8'hC0; 15'h0237: d <= 8'hC0;
                15'h0238: d <= 8'hC0; 15'h0239: d <= 8'hC0; 15'h023A: d <= 8'hC0; 15'h023B: d <= 8'hC0;
                15'h023C: d <= 8'hC0; 15'h023D: d <= 8'hC0; 15'h023E: d <= 8'hC0; 15'h023F: d <= 8'hC0;
                15'h0240: d <= 8'hC0; 15'h0241: d <= 8'hC0; 15'h0242: d <= 8'hC0; 15'h0243: d <= 8'hC0;
                15'h0244: d <= 8'hC0; 15'h0245: d <= 8'hC0; 15'h0246: d <= 8'hC0; 15'h0247: d <= 8'hC0;
                15'h0248: d <= 8'hC0; 15'h0249: d <= 8'hC0; 15'h024A: d <= 8'hC0; 15'h024B: d <= 8'hC0;
                15'h024C: d <= 8'hC0; 15'h024D: d <= 8'hC0; 15'h024E: d <= 8'hC0; 15'h024F: d <= 8'hC0;
                15'h0250: d <= 8'hC0; 15'h0251: d <= 8'hC0; 15'h0252: d <= 8'hC0; 15'h0253: d <= 8'hC0;
                15'h0254: d <= 8'hC0; 15'h0255: d <= 8'hC0; 15'h0256: d <= 8'hC0; 15'h0257: d <= 8'hC0;
                15'h0258: d <= 8'hC0; 15'h0259: d <= 8'hC0; 15'h025A: d <= 8'hC0; 15'h025B: d <= 8'hC0;
                15'h025C: d <= 8'hC0; 15'h025D: d <= 8'hC0; 15'h025E: d <= 8'hC0; 15'h025F: d <= 8'hC0;
                15'h0260: d <= 8'hC0; 15'h0261: d <= 8'hC0; 15'h0262: d <= 8'hC0; 15'h0263: d <= 8'hC0;
                15'h0264: d <= 8'hC0; 15'h0265: d <= 8'hC0; 15'h0266: d <= 8'hC0; 15'h0267: d <= 8'hC0;
                15'h0268: d <= 8'hC0; 15'h0269: d <= 8'hC0; 15'h026A: d <= 8'hC0; 15'h026B: d <= 8'hC0;
                15'h026C: d <= 8'hC0; 15'h026D: d <= 8'hC0; 15'h026E: d <= 8'hC0; 15'h026F: d <= 8'hC0;
                15'h0270: d <= 8'hC0; 15'h0271: d <= 8'hC0; 15'h0272: d <= 8'hC0; 15'h0273: d <= 8'hC0;
                15'h0274: d <= 8'hC0; 15'h0275: d <= 8'hC0; 15'h0276: d <= 8'hC0; 15'h0277: d <= 8'hC0;
                15'h0278: d <= 8'hC0; 15'h0279: d <= 8'hC0; 15'h027A: d <= 8'hC0; 15'h027B: d <= 8'hC0;
                15'h027C: d <= 8'hC0; 15'h027D: d <= 8'hC0; 15'h027E: d <= 8'hC0; 15'h027F: d <= 8'hC0;
                15'h0280: d <= 8'hC0; 15'h0281: d <= 8'hC0; 15'h0282: d <= 8'hC0; 15'h0283: d <= 8'hC0;
                15'h0284: d <= 8'hC0; 15'h0285: d <= 8'hC0; 15'h0286: d <= 8'hC0; 15'h0287: d <= 8'hC0;
                15'h0288: d <= 8'hC0; 15'h0289: d <= 8'hC0; 15'h028A: d <= 8'hC0; 15'h028B: d <= 8'hC0;
                15'h028C: d <= 8'hC0; 15'h028D: d <= 8'hC0; 15'h028E: d <= 8'hC0; 15'h028F: d <= 8'hC0;
                15'h0290: d <= 8'hC0; 15'h0291: d <= 8'hC0; 15'h0292: d <= 8'hC0; 15'h0293: d <= 8'hC0;
                15'h0294: d <= 8'hC0; 15'h0295: d <= 8'hC0; 15'h0296: d <= 8'hC0; 15'h0297: d <= 8'hC0;
                15'h0298: d <= 8'hC0; 15'h0299: d <= 8'hC0; 15'h029A: d <= 8'hC0; 15'h029B: d <= 8'hC0;
                15'h029C: d <= 8'hC0; 15'h029D: d <= 8'hC0; 15'h029E: d <= 8'hC0; 15'h029F: d <= 8'hC0;
                15'h02A0: d <= 8'hC0; 15'h02A1: d <= 8'hC0; 15'h02A2: d <= 8'hC0; 15'h02A3: d <= 8'hC0;
                15'h02A4: d <= 8'hC0; 15'h02A5: d <= 8'hC0; 15'h02A6: d <= 8'hC0; 15'h02A7: d <= 8'hC0;
                15'h02A8: d <= 8'hC0; 15'h02A9: d <= 8'hC0; 15'h02AA: d <= 8'hC0; 15'h02AB: d <= 8'hC0;
                15'h02AC: d <= 8'hC0; 15'h02AD: d <= 8'hC0; 15'h02AE: d <= 8'hC0; 15'h02AF: d <= 8'hC0;
                15'h02B0: d <= 8'hC0; 15'h02B1: d <= 8'hC0; 15'h02B2: d <= 8'hC0; 15'h02B3: d <= 8'hC0;
                15'h02B4: d <= 8'hC0; 15'h02B5: d <= 8'hC0; 15'h02B6: d <= 8'hC0; 15'h02B7: d <= 8'hC0;
                15'h02B8: d <= 8'hC0; 15'h02B9: d <= 8'hC0; 15'h02BA: d <= 8'hC0; 15'h02BB: d <= 8'hC0;
                15'h02BC: d <= 8'hC0; 15'h02BD: d <= 8'hC0; 15'h02BE: d <= 8'hC0; 15'h02BF: d <= 8'hC0;
                15'h02C0: d <= 8'hC0; 15'h02C1: d <= 8'hC0; 15'h02C2: d <= 8'hC0; 15'h02C3: d <= 8'hC0;
                15'h02C4: d <= 8'hC0; 15'h02C5: d <= 8'hC0; 15'h02C6: d <= 8'hC0; 15'h02C7: d <= 8'hC0;
                15'h02C8: d <= 8'hC0; 15'h02C9: d <= 8'hC0; 15'h02CA: d <= 8'hC0; 15'h02CB: d <= 8'hC0;
                15'h02CC: d <= 8'hC0; 15'h02CD: d <= 8'hC0; 15'h02CE: d <= 8'hC0; 15'h02CF: d <= 8'hC0;
                15'h02D0: d <= 8'hC0; 15'h02D1: d <= 8'hC0; 15'h02D2: d <= 8'hC0; 15'h02D3: d <= 8'hC0;
                15'h02D4: d <= 8'hC0; 15'h02D5: d <= 8'hC0; 15'h02D6: d <= 8'hC0; 15'h02D7: d <= 8'hC0;
                15'h02D8: d <= 8'hC0; 15'h02D9: d <= 8'hC0; 15'h02DA: d <= 8'hC0; 15'h02DB: d <= 8'hC0;
                15'h02DC: d <= 8'hC0; 15'h02DD: d <= 8'hC0; 15'h02DE: d <= 8'hC0; 15'h02DF: d <= 8'hC0;
                15'h02E0: d <= 8'hC0; 15'h02E1: d <= 8'hC0; 15'h02E2: d <= 8'hC0; 15'h02E3: d <= 8'hC0;
                15'h02E4: d <= 8'hC0; 15'h02E5: d <= 8'hC0; 15'h02E6: d <= 8'hC0; 15'h02E7: d <= 8'hC0;
                15'h02E8: d <= 8'hC0; 15'h02E9: d <= 8'hC0; 15'h02EA: d <= 8'hC0; 15'h02EB: d <= 8'hC0;
                15'h02EC: d <= 8'hC0; 15'h02ED: d <= 8'hC0; 15'h02EE: d <= 8'hC0; 15'h02EF: d <= 8'hC0;
                15'h02F0: d <= 8'hC0; 15'h02F1: d <= 8'hC0; 15'h02F2: d <= 8'hC0; 15'h02F3: d <= 8'hC0;
                15'h02F4: d <= 8'hC0; 15'h02F5: d <= 8'hC0; 15'h02F6: d <= 8'hC0; 15'h02F7: d <= 8'hC0;
                15'h02F8: d <= 8'hC0; 15'h02F9: d <= 8'hC0; 15'h02FA: d <= 8'hC0; 15'h02FB: d <= 8'hC0;
                15'h02FC: d <= 8'hC0; 15'h02FD: d <= 8'hC0; 15'h02FE: d <= 8'hC0; 15'h02FF: d <= 8'hC0;
                15'h0300: d <= 8'hC0; 15'h0301: d <= 8'hC0; 15'h0302: d <= 8'hC0; 15'h0303: d <= 8'hC0;
                15'h0304: d <= 8'hC0; 15'h0305: d <= 8'hC0; 15'h0306: d <= 8'hC0; 15'h0307: d <= 8'hC0;
                15'h0308: d <= 8'hC0; 15'h0309: d <= 8'hC0; 15'h030A: d <= 8'hC0; 15'h030B: d <= 8'hC0;
                15'h030C: d <= 8'hC0; 15'h030D: d <= 8'hC0; 15'h030E: d <= 8'hC0; 15'h030F: d <= 8'hC0;
                15'h0310: d <= 8'hC0; 15'h0311: d <= 8'hC0; 15'h0312: d <= 8'hC0; 15'h0313: d <= 8'hC0;
                15'h0314: d <= 8'hC0; 15'h0315: d <= 8'hC0; 15'h0316: d <= 8'hC0; 15'h0317: d <= 8'hC0;
                15'h0318: d <= 8'hC0; 15'h0319: d <= 8'hC0; 15'h031A: d <= 8'hC0; 15'h031B: d <= 8'hC0;
                15'h031C: d <= 8'hC0; 15'h031D: d <= 8'hC0; 15'h031E: d <= 8'hC0; 15'h031F: d <= 8'hC0;
                15'h0320: d <= 8'hC0; 15'h0321: d <= 8'hC0; 15'h0322: d <= 8'hC0; 15'h0323: d <= 8'hC0;
                15'h0324: d <= 8'hC0; 15'h0325: d <= 8'hC0; 15'h0326: d <= 8'hC0; 15'h0327: d <= 8'hC0;
                15'h0328: d <= 8'hC0; 15'h0329: d <= 8'hC0; 15'h032A: d <= 8'hC0; 15'h032B: d <= 8'hC0;
                15'h032C: d <= 8'hC0; 15'h032D: d <= 8'hC0; 15'h032E: d <= 8'hC0; 15'h032F: d <= 8'hC0;
                15'h0330: d <= 8'hC0; 15'h0331: d <= 8'hC0; 15'h0332: d <= 8'hC0; 15'h0333: d <= 8'hC0;
                15'h0334: d <= 8'hC0; 15'h0335: d <= 8'hC0; 15'h0336: d <= 8'hC0; 15'h0337: d <= 8'hC0;
                15'h0338: d <= 8'hC0; 15'h0339: d <= 8'hC0; 15'h033A: d <= 8'hC0; 15'h033B: d <= 8'hC0;
                15'h033C: d <= 8'hC0; 15'h033D: d <= 8'hC0; 15'h033E: d <= 8'hC0; 15'h033F: d <= 8'hC0;
                15'h0340: d <= 8'hC0; 15'h0341: d <= 8'hC0; 15'h0342: d <= 8'hC0; 15'h0343: d <= 8'hC0;
                15'h0344: d <= 8'hC0; 15'h0345: d <= 8'hC0; 15'h0346: d <= 8'hC0; 15'h0347: d <= 8'hC0;
                15'h0348: d <= 8'hC0; 15'h0349: d <= 8'hC0; 15'h034A: d <= 8'hC0; 15'h034B: d <= 8'hC0;
                15'h034C: d <= 8'hC0; 15'h034D: d <= 8'hC0; 15'h034E: d <= 8'hC0; 15'h034F: d <= 8'hC0;
                15'h0350: d <= 8'hC0; 15'h0351: d <= 8'hC0; 15'h0352: d <= 8'hC0; 15'h0353: d <= 8'hC0;
                15'h0354: d <= 8'hC0; 15'h0355: d <= 8'hC0; 15'h0356: d <= 8'hC0; 15'h0357: d <= 8'hC0;
                15'h0358: d <= 8'hC0; 15'h0359: d <= 8'hC0; 15'h035A: d <= 8'hC0; 15'h035B: d <= 8'hC0;
                15'h035C: d <= 8'hC0; 15'h035D: d <= 8'hC0; 15'h035E: d <= 8'hC0; 15'h035F: d <= 8'hC0;
                15'h0360: d <= 8'hC0; 15'h0361: d <= 8'hC0; 15'h0362: d <= 8'hC0; 15'h0363: d <= 8'hC0;
                15'h0364: d <= 8'hC0; 15'h0365: d <= 8'hC0; 15'h0366: d <= 8'hC0; 15'h0367: d <= 8'hC0;
                15'h0368: d <= 8'hC0; 15'h0369: d <= 8'hC0; 15'h036A: d <= 8'hC0; 15'h036B: d <= 8'hC0;
                15'h036C: d <= 8'hC0; 15'h036D: d <= 8'hC0; 15'h036E: d <= 8'hC0; 15'h036F: d <= 8'hC0;
                15'h0370: d <= 8'hC0; 15'h0371: d <= 8'hC0; 15'h0372: d <= 8'hC0; 15'h0373: d <= 8'hC0;
                15'h0374: d <= 8'hC0; 15'h0375: d <= 8'hC0; 15'h0376: d <= 8'hC0; 15'h0377: d <= 8'hC0;
                15'h0378: d <= 8'hC0; 15'h0379: d <= 8'hC0; 15'h037A: d <= 8'hC0; 15'h037B: d <= 8'hC0;
                15'h037C: d <= 8'hC0; 15'h037D: d <= 8'hC0; 15'h037E: d <= 8'hC0; 15'h037F: d <= 8'hC0;
                15'h0380: d <= 8'hC0; 15'h0381: d <= 8'hC0; 15'h0382: d <= 8'hC0; 15'h0383: d <= 8'hC0;
                15'h0384: d <= 8'hC0; 15'h0385: d <= 8'hC0; 15'h0386: d <= 8'hC0; 15'h0387: d <= 8'hC0;
                15'h0388: d <= 8'hC0; 15'h0389: d <= 8'hC0; 15'h038A: d <= 8'hC0; 15'h038B: d <= 8'hC0;
                15'h038C: d <= 8'hC0; 15'h038D: d <= 8'hC0; 15'h038E: d <= 8'hC0; 15'h038F: d <= 8'hC0;
                15'h0390: d <= 8'hC0; 15'h0391: d <= 8'hC0; 15'h0392: d <= 8'hC0; 15'h0393: d <= 8'hC0;
                15'h0394: d <= 8'hC0; 15'h0395: d <= 8'hC0; 15'h0396: d <= 8'hC0; 15'h0397: d <= 8'hC0;
                15'h0398: d <= 8'hC0; 15'h0399: d <= 8'hC0; 15'h039A: d <= 8'hC0; 15'h039B: d <= 8'hC0;
                15'h039C: d <= 8'hC0; 15'h039D: d <= 8'hC0; 15'h039E: d <= 8'hC0; 15'h039F: d <= 8'hC0;
                15'h03A0: d <= 8'hC0; 15'h03A1: d <= 8'hC0; 15'h03A2: d <= 8'hC0; 15'h03A3: d <= 8'hC0;
                15'h03A4: d <= 8'hC0; 15'h03A5: d <= 8'hC0; 15'h03A6: d <= 8'hC0; 15'h03A7: d <= 8'hC0;
                15'h03A8: d <= 8'hC0; 15'h03A9: d <= 8'hC0; 15'h03AA: d <= 8'hC0; 15'h03AB: d <= 8'hC0;
                15'h03AC: d <= 8'hC0; 15'h03AD: d <= 8'hC0; 15'h03AE: d <= 8'hC0; 15'h03AF: d <= 8'hC0;
                15'h03B0: d <= 8'hC0; 15'h03B1: d <= 8'hC0; 15'h03B2: d <= 8'hC0; 15'h03B3: d <= 8'hC0;
                15'h03B4: d <= 8'hC0; 15'h03B5: d <= 8'hC0; 15'h03B6: d <= 8'hC0; 15'h03B7: d <= 8'hC0;
                15'h03B8: d <= 8'hC0; 15'h03B9: d <= 8'hC0; 15'h03BA: d <= 8'hC0; 15'h03BB: d <= 8'hC0;
                15'h03BC: d <= 8'hC0; 15'h03BD: d <= 8'hC0; 15'h03BE: d <= 8'hC0; 15'h03BF: d <= 8'hC0;
                15'h03C0: d <= 8'hC0; 15'h03C1: d <= 8'hC0; 15'h03C2: d <= 8'hC0; 15'h03C3: d <= 8'hC0;
                15'h03C4: d <= 8'hC0; 15'h03C5: d <= 8'hC0; 15'h03C6: d <= 8'hC0; 15'h03C7: d <= 8'hC0;
                15'h03C8: d <= 8'hC0; 15'h03C9: d <= 8'hC0; 15'h03CA: d <= 8'hC0; 15'h03CB: d <= 8'hC0;
                15'h03CC: d <= 8'hC0; 15'h03CD: d <= 8'hC0; 15'h03CE: d <= 8'hC0; 15'h03CF: d <= 8'hC0;
                15'h03D0: d <= 8'hC0; 15'h03D1: d <= 8'hC0; 15'h03D2: d <= 8'hC0; 15'h03D3: d <= 8'hC0;
                15'h03D4: d <= 8'hC0; 15'h03D5: d <= 8'hC0; 15'h03D6: d <= 8'hC0; 15'h03D7: d <= 8'hC0;
                15'h03D8: d <= 8'hC0; 15'h03D9: d <= 8'hC0; 15'h03DA: d <= 8'hC0; 15'h03DB: d <= 8'hC0;
                15'h03DC: d <= 8'hC0; 15'h03DD: d <= 8'hC0; 15'h03DE: d <= 8'hC0; 15'h03DF: d <= 8'hC0;
                15'h03E0: d <= 8'hC0; 15'h03E1: d <= 8'hC0; 15'h03E2: d <= 8'hC0; 15'h03E3: d <= 8'hC0;
                15'h03E4: d <= 8'hC0; 15'h03E5: d <= 8'hC0; 15'h03E6: d <= 8'hC0; 15'h03E7: d <= 8'hC0;
                15'h03E8: d <= 8'hC0; 15'h03E9: d <= 8'hC0; 15'h03EA: d <= 8'hC0; 15'h03EB: d <= 8'hC0;
                15'h03EC: d <= 8'hC0; 15'h03ED: d <= 8'hC0; 15'h03EE: d <= 8'hC0; 15'h03EF: d <= 8'hC0;
                15'h03F0: d <= 8'hC0; 15'h03F1: d <= 8'hC0; 15'h03F2: d <= 8'hC0; 15'h03F3: d <= 8'hC0;
                15'h03F4: d <= 8'hC0; 15'h03F5: d <= 8'hC0; 15'h03F6: d <= 8'hC0; 15'h03F7: d <= 8'hC0;
                15'h03F8: d <= 8'hC0; 15'h03F9: d <= 8'hC0; 15'h03FA: d <= 8'hC0; 15'h03FB: d <= 8'hC0;
                15'h03FC: d <= 8'hC0; 15'h03FD: d <= 8'hC0; 15'h03FE: d <= 8'hC0; 15'h03FF: d <= 8'hC0;
                15'h0400: d <= 8'hC0; 15'h0401: d <= 8'hC0; 15'h0402: d <= 8'hC0; 15'h0403: d <= 8'hC0;
                15'h0404: d <= 8'hC0; 15'h0405: d <= 8'hC0; 15'h0406: d <= 8'hC0; 15'h0407: d <= 8'hC0;
                15'h0408: d <= 8'hC0; 15'h0409: d <= 8'hC0; 15'h040A: d <= 8'hC0; 15'h040B: d <= 8'hC0;
                15'h040C: d <= 8'hC0; 15'h040D: d <= 8'hC0; 15'h040E: d <= 8'hC0; 15'h040F: d <= 8'hC0;
                15'h0410: d <= 8'hC0; 15'h0411: d <= 8'hC0; 15'h0412: d <= 8'hC0; 15'h0413: d <= 8'hC0;
                15'h0414: d <= 8'hC0; 15'h0415: d <= 8'hC0; 15'h0416: d <= 8'hC0; 15'h0417: d <= 8'hC0;
                15'h0418: d <= 8'hC0; 15'h0419: d <= 8'hC0; 15'h041A: d <= 8'hC0; 15'h041B: d <= 8'hC0;
                15'h041C: d <= 8'hC0; 15'h041D: d <= 8'hC0; 15'h041E: d <= 8'hC0; 15'h041F: d <= 8'hC0;
                15'h0420: d <= 8'hC0; 15'h0421: d <= 8'hC0; 15'h0422: d <= 8'hC0; 15'h0423: d <= 8'hC0;
                15'h0424: d <= 8'hC0; 15'h0425: d <= 8'hC0; 15'h0426: d <= 8'hC0; 15'h0427: d <= 8'hC0;
                15'h0428: d <= 8'hC0; 15'h0429: d <= 8'hC0; 15'h042A: d <= 8'hC0; 15'h042B: d <= 8'hC0;
                15'h042C: d <= 8'hC0; 15'h042D: d <= 8'hC0; 15'h042E: d <= 8'hC0; 15'h042F: d <= 8'hC0;
                15'h0430: d <= 8'hC0; 15'h0431: d <= 8'hC0; 15'h0432: d <= 8'hC0; 15'h0433: d <= 8'hC0;
                15'h0434: d <= 8'hC0; 15'h0435: d <= 8'hC0; 15'h0436: d <= 8'hC0; 15'h0437: d <= 8'hC0;
                15'h0438: d <= 8'hC0; 15'h0439: d <= 8'hC0; 15'h043A: d <= 8'hC0; 15'h043B: d <= 8'hC0;
                15'h043C: d <= 8'hC0; 15'h043D: d <= 8'hC0; 15'h043E: d <= 8'hC0; 15'h043F: d <= 8'hC0;
                15'h0440: d <= 8'hC0; 15'h0441: d <= 8'hC0; 15'h0442: d <= 8'hC0; 15'h0443: d <= 8'hC0;
                15'h0444: d <= 8'hC0; 15'h0445: d <= 8'hC0; 15'h0446: d <= 8'hC0; 15'h0447: d <= 8'hC0;
                15'h0448: d <= 8'hC0; 15'h0449: d <= 8'hC0; 15'h044A: d <= 8'hC0; 15'h044B: d <= 8'hC0;
                15'h044C: d <= 8'hC0; 15'h044D: d <= 8'hC0; 15'h044E: d <= 8'hC0; 15'h044F: d <= 8'hC0;
                15'h0450: d <= 8'hC0; 15'h0451: d <= 8'hC0; 15'h0452: d <= 8'hC0; 15'h0453: d <= 8'hC0;
                15'h0454: d <= 8'hC0; 15'h0455: d <= 8'hC0; 15'h0456: d <= 8'hC0; 15'h0457: d <= 8'hC0;
                15'h0458: d <= 8'hC0; 15'h0459: d <= 8'hC0; 15'h045A: d <= 8'hC0; 15'h045B: d <= 8'hC0;
                15'h045C: d <= 8'hC0; 15'h045D: d <= 8'hC0; 15'h045E: d <= 8'hC0; 15'h045F: d <= 8'hC0;
                15'h0460: d <= 8'hC0; 15'h0461: d <= 8'hC0; 15'h0462: d <= 8'hC0; 15'h0463: d <= 8'hC0;
                15'h0464: d <= 8'hC0; 15'h0465: d <= 8'hC0; 15'h0466: d <= 8'hC0; 15'h0467: d <= 8'hC0;
                15'h0468: d <= 8'hC0; 15'h0469: d <= 8'hC0; 15'h046A: d <= 8'hC0; 15'h046B: d <= 8'hC0;
                15'h046C: d <= 8'hC0; 15'h046D: d <= 8'hC0; 15'h046E: d <= 8'hC0; 15'h046F: d <= 8'hC0;
                15'h0470: d <= 8'hC0; 15'h0471: d <= 8'hC0; 15'h0472: d <= 8'hC0; 15'h0473: d <= 8'hC0;
                15'h0474: d <= 8'hC0; 15'h0475: d <= 8'hC0; 15'h0476: d <= 8'hC0; 15'h0477: d <= 8'hC0;
                15'h0478: d <= 8'hC0; 15'h0479: d <= 8'hC0; 15'h047A: d <= 8'hC0; 15'h047B: d <= 8'hC0;
                15'h047C: d <= 8'hC0; 15'h047D: d <= 8'hC0; 15'h047E: d <= 8'hC0; 15'h047F: d <= 8'hC0;
                15'h0480: d <= 8'hC0; 15'h0481: d <= 8'hC0; 15'h0482: d <= 8'hC0; 15'h0483: d <= 8'hC0;
                15'h0484: d <= 8'hC0; 15'h0485: d <= 8'hC0; 15'h0486: d <= 8'hC0; 15'h0487: d <= 8'hC0;
                15'h0488: d <= 8'hC0; 15'h0489: d <= 8'hC0; 15'h048A: d <= 8'hC0; 15'h048B: d <= 8'hC0;
                15'h048C: d <= 8'hC0; 15'h048D: d <= 8'hC0; 15'h048E: d <= 8'hC0; 15'h048F: d <= 8'hC0;
                15'h0490: d <= 8'hC0; 15'h0491: d <= 8'hC0; 15'h0492: d <= 8'hC0; 15'h0493: d <= 8'hC0;
                15'h0494: d <= 8'hC0; 15'h0495: d <= 8'hC0; 15'h0496: d <= 8'hC0; 15'h0497: d <= 8'hC0;
                15'h0498: d <= 8'hC0; 15'h0499: d <= 8'hC0; 15'h049A: d <= 8'hC0; 15'h049B: d <= 8'hC0;
                15'h049C: d <= 8'hC0; 15'h049D: d <= 8'hC0; 15'h049E: d <= 8'hC0; 15'h049F: d <= 8'hC0;
                15'h04A0: d <= 8'hC0; 15'h04A1: d <= 8'hC0; 15'h04A2: d <= 8'hC0; 15'h04A3: d <= 8'hC0;
                15'h04A4: d <= 8'hC0; 15'h04A5: d <= 8'hC0; 15'h04A6: d <= 8'hC0; 15'h04A7: d <= 8'hC0;
                15'h04A8: d <= 8'hC0; 15'h04A9: d <= 8'hC0; 15'h04AA: d <= 8'hC0; 15'h04AB: d <= 8'hC0;
                15'h04AC: d <= 8'hC0; 15'h04AD: d <= 8'hC0; 15'h04AE: d <= 8'hC0; 15'h04AF: d <= 8'hC0;
                15'h04B0: d <= 8'hC0; 15'h04B1: d <= 8'hC0; 15'h04B2: d <= 8'hC0; 15'h04B3: d <= 8'hC0;
                15'h04B4: d <= 8'hC0; 15'h04B5: d <= 8'hC0; 15'h04B6: d <= 8'hC0; 15'h04B7: d <= 8'hC0;
                15'h04B8: d <= 8'hC0; 15'h04B9: d <= 8'hC0; 15'h04BA: d <= 8'hC0; 15'h04BB: d <= 8'hC0;
                15'h04BC: d <= 8'hC0; 15'h04BD: d <= 8'hC0; 15'h04BE: d <= 8'hC0; 15'h04BF: d <= 8'hC0;
                15'h04C0: d <= 8'hC0; 15'h04C1: d <= 8'hC0; 15'h04C2: d <= 8'hC0; 15'h04C3: d <= 8'hC0;
                15'h04C4: d <= 8'hC0; 15'h04C5: d <= 8'hC0; 15'h04C6: d <= 8'hC0; 15'h04C7: d <= 8'hC0;
                15'h04C8: d <= 8'hC0; 15'h04C9: d <= 8'hC0; 15'h04CA: d <= 8'hC0; 15'h04CB: d <= 8'hC0;
                15'h04CC: d <= 8'hC0; 15'h04CD: d <= 8'hC0; 15'h04CE: d <= 8'hC0; 15'h04CF: d <= 8'hC0;
                15'h04D0: d <= 8'hC0; 15'h04D1: d <= 8'hC0; 15'h04D2: d <= 8'hC0; 15'h04D3: d <= 8'hC0;
                15'h04D4: d <= 8'hC0; 15'h04D5: d <= 8'hC0; 15'h04D6: d <= 8'hC0; 15'h04D7: d <= 8'hC0;
                15'h04D8: d <= 8'hC0; 15'h04D9: d <= 8'hC0; 15'h04DA: d <= 8'hC0; 15'h04DB: d <= 8'hC0;
                15'h04DC: d <= 8'hC0; 15'h04DD: d <= 8'hC0; 15'h04DE: d <= 8'hC0; 15'h04DF: d <= 8'hC0;
                15'h04E0: d <= 8'hC0; 15'h04E1: d <= 8'hC0; 15'h04E2: d <= 8'hC0; 15'h04E3: d <= 8'hC0;
                15'h04E4: d <= 8'hC0; 15'h04E5: d <= 8'hC0; 15'h04E6: d <= 8'hC0; 15'h04E7: d <= 8'hC0;
                15'h04E8: d <= 8'hC0; 15'h04E9: d <= 8'hC0; 15'h04EA: d <= 8'hC0; 15'h04EB: d <= 8'hC0;
                15'h04EC: d <= 8'hC0; 15'h04ED: d <= 8'hC0; 15'h04EE: d <= 8'hC0; 15'h04EF: d <= 8'hC0;
                15'h04F0: d <= 8'hC0; 15'h04F1: d <= 8'hC0; 15'h04F2: d <= 8'hC0; 15'h04F3: d <= 8'hC0;
                15'h04F4: d <= 8'hC0; 15'h04F5: d <= 8'hC0; 15'h04F6: d <= 8'hC0; 15'h04F7: d <= 8'hC0;
                15'h04F8: d <= 8'hC0; 15'h04F9: d <= 8'hC0; 15'h04FA: d <= 8'hC0; 15'h04FB: d <= 8'hC0;
                15'h04FC: d <= 8'hC0; 15'h04FD: d <= 8'hC0; 15'h04FE: d <= 8'hC0; 15'h04FF: d <= 8'hC0;
                15'h0500: d <= 8'hC0; 15'h0501: d <= 8'hC0; 15'h0502: d <= 8'hC0; 15'h0503: d <= 8'hC0;
                15'h0504: d <= 8'hC0; 15'h0505: d <= 8'hC0; 15'h0506: d <= 8'hC0; 15'h0507: d <= 8'hC0;
                15'h0508: d <= 8'hC0; 15'h0509: d <= 8'hC0; 15'h050A: d <= 8'hC0; 15'h050B: d <= 8'hC0;
                15'h050C: d <= 8'hC0; 15'h050D: d <= 8'hC0; 15'h050E: d <= 8'hC0; 15'h050F: d <= 8'hC0;
                15'h0510: d <= 8'hC0; 15'h0511: d <= 8'hC0; 15'h0512: d <= 8'hC0; 15'h0513: d <= 8'hC0;
                15'h0514: d <= 8'hC0; 15'h0515: d <= 8'hC0; 15'h0516: d <= 8'hC0; 15'h0517: d <= 8'hC0;
                15'h0518: d <= 8'hC0; 15'h0519: d <= 8'hC0; 15'h051A: d <= 8'hC0; 15'h051B: d <= 8'hC0;
                15'h051C: d <= 8'hC0; 15'h051D: d <= 8'hC0; 15'h051E: d <= 8'hC0; 15'h051F: d <= 8'hC0;
                15'h0520: d <= 8'hC0; 15'h0521: d <= 8'hC0; 15'h0522: d <= 8'hC0; 15'h0523: d <= 8'hC0;
                15'h0524: d <= 8'hC0; 15'h0525: d <= 8'hC0; 15'h0526: d <= 8'hC0; 15'h0527: d <= 8'hC0;
                15'h0528: d <= 8'hC0; 15'h0529: d <= 8'hC0; 15'h052A: d <= 8'hC0; 15'h052B: d <= 8'hC0;
                15'h052C: d <= 8'hC0; 15'h052D: d <= 8'hC0; 15'h052E: d <= 8'hC0; 15'h052F: d <= 8'hC0;
                15'h0530: d <= 8'hC0; 15'h0531: d <= 8'hC0; 15'h0532: d <= 8'hC0; 15'h0533: d <= 8'hC0;
                15'h0534: d <= 8'hC0; 15'h0535: d <= 8'hC0; 15'h0536: d <= 8'hC0; 15'h0537: d <= 8'hC0;
                15'h0538: d <= 8'hC0; 15'h0539: d <= 8'hC0; 15'h053A: d <= 8'hC0; 15'h053B: d <= 8'hC0;
                15'h053C: d <= 8'hC0; 15'h053D: d <= 8'hC0; 15'h053E: d <= 8'hC0; 15'h053F: d <= 8'hC0;
                15'h0540: d <= 8'hC0; 15'h0541: d <= 8'hC0; 15'h0542: d <= 8'hC0; 15'h0543: d <= 8'hC0;
                15'h0544: d <= 8'hC0; 15'h0545: d <= 8'hC0; 15'h0546: d <= 8'hC0; 15'h0547: d <= 8'hC0;
                15'h0548: d <= 8'hC0; 15'h0549: d <= 8'hC0; 15'h054A: d <= 8'hC0; 15'h054B: d <= 8'hC0;
                15'h054C: d <= 8'hC0; 15'h054D: d <= 8'hC0; 15'h054E: d <= 8'hC0; 15'h054F: d <= 8'hC0;
                15'h0550: d <= 8'hC0; 15'h0551: d <= 8'hC0; 15'h0552: d <= 8'hC0; 15'h0553: d <= 8'hC0;
                15'h0554: d <= 8'hC0; 15'h0555: d <= 8'hC0; 15'h0556: d <= 8'hC0; 15'h0557: d <= 8'hC0;
                15'h0558: d <= 8'hC0; 15'h0559: d <= 8'hC0; 15'h055A: d <= 8'hC0; 15'h055B: d <= 8'hC0;
                15'h055C: d <= 8'hC0; 15'h055D: d <= 8'hC0; 15'h055E: d <= 8'hC0; 15'h055F: d <= 8'hC0;
                15'h0560: d <= 8'hC0; 15'h0561: d <= 8'hC0; 15'h0562: d <= 8'hC0; 15'h0563: d <= 8'hC0;
                15'h0564: d <= 8'hC0; 15'h0565: d <= 8'hC0; 15'h0566: d <= 8'hC0; 15'h0567: d <= 8'hC0;
                15'h0568: d <= 8'hC0; 15'h0569: d <= 8'hC0; 15'h056A: d <= 8'hC0; 15'h056B: d <= 8'hC0;
                15'h056C: d <= 8'hC0; 15'h056D: d <= 8'hC0; 15'h056E: d <= 8'hC0; 15'h056F: d <= 8'hC0;
                15'h0570: d <= 8'hC0; 15'h0571: d <= 8'hC0; 15'h0572: d <= 8'hC0; 15'h0573: d <= 8'hC0;
                15'h0574: d <= 8'hC0; 15'h0575: d <= 8'hC0; 15'h0576: d <= 8'hC0; 15'h0577: d <= 8'hC0;
                15'h0578: d <= 8'hC0; 15'h0579: d <= 8'hC0; 15'h057A: d <= 8'hC0; 15'h057B: d <= 8'hC0;
                15'h057C: d <= 8'hC0; 15'h057D: d <= 8'hC0; 15'h057E: d <= 8'hC0; 15'h057F: d <= 8'hC0;
                15'h0580: d <= 8'hC0; 15'h0581: d <= 8'hC0; 15'h0582: d <= 8'hC0; 15'h0583: d <= 8'hC0;
                15'h0584: d <= 8'hC0; 15'h0585: d <= 8'hC0; 15'h0586: d <= 8'hC0; 15'h0587: d <= 8'hC0;
                15'h0588: d <= 8'hC0; 15'h0589: d <= 8'hC0; 15'h058A: d <= 8'hC0; 15'h058B: d <= 8'hC0;
                15'h058C: d <= 8'hC0; 15'h058D: d <= 8'hC0; 15'h058E: d <= 8'hC0; 15'h058F: d <= 8'hC0;
                15'h0590: d <= 8'hC0; 15'h0591: d <= 8'hC0; 15'h0592: d <= 8'hC0; 15'h0593: d <= 8'hC0;
                15'h0594: d <= 8'hC0; 15'h0595: d <= 8'hC0; 15'h0596: d <= 8'hC0; 15'h0597: d <= 8'hC0;
                15'h0598: d <= 8'hC0; 15'h0599: d <= 8'hC0; 15'h059A: d <= 8'hC0; 15'h059B: d <= 8'hC0;
                15'h059C: d <= 8'hC0; 15'h059D: d <= 8'hC0; 15'h059E: d <= 8'hC0; 15'h059F: d <= 8'hC0;
                15'h05A0: d <= 8'hC0; 15'h05A1: d <= 8'hC0; 15'h05A2: d <= 8'hC0; 15'h05A3: d <= 8'hC0;
                15'h05A4: d <= 8'hC0; 15'h05A5: d <= 8'hC0; 15'h05A6: d <= 8'hC0; 15'h05A7: d <= 8'hC0;
                15'h05A8: d <= 8'hC0; 15'h05A9: d <= 8'hC0; 15'h05AA: d <= 8'hC0; 15'h05AB: d <= 8'hC0;
                15'h05AC: d <= 8'hC0; 15'h05AD: d <= 8'hC0; 15'h05AE: d <= 8'hC0; 15'h05AF: d <= 8'hC0;
                15'h05B0: d <= 8'hC0; 15'h05B1: d <= 8'hC0; 15'h05B2: d <= 8'hC0; 15'h05B3: d <= 8'hC0;
                15'h05B4: d <= 8'hC0; 15'h05B5: d <= 8'hC0; 15'h05B6: d <= 8'hC0; 15'h05B7: d <= 8'hC0;
                15'h05B8: d <= 8'hC0; 15'h05B9: d <= 8'hC0; 15'h05BA: d <= 8'hC0; 15'h05BB: d <= 8'hC0;
                15'h05BC: d <= 8'hC0; 15'h05BD: d <= 8'hC0; 15'h05BE: d <= 8'hC0; 15'h05BF: d <= 8'hC0;
                15'h05C0: d <= 8'hC0; 15'h05C1: d <= 8'hC0; 15'h05C2: d <= 8'hC0; 15'h05C3: d <= 8'hC0;
                15'h05C4: d <= 8'hC0; 15'h05C5: d <= 8'hC0; 15'h05C6: d <= 8'hC0; 15'h05C7: d <= 8'hC0;
                15'h05C8: d <= 8'hC0; 15'h05C9: d <= 8'hC0; 15'h05CA: d <= 8'hC0; 15'h05CB: d <= 8'hC0;
                15'h05CC: d <= 8'hC0; 15'h05CD: d <= 8'hC0; 15'h05CE: d <= 8'hC0; 15'h05CF: d <= 8'hC0;
                15'h05D0: d <= 8'hC0; 15'h05D1: d <= 8'hC0; 15'h05D2: d <= 8'hC0; 15'h05D3: d <= 8'hC0;
                15'h05D4: d <= 8'hC0; 15'h05D5: d <= 8'hC0; 15'h05D6: d <= 8'hC0; 15'h05D7: d <= 8'hC0;
                15'h05D8: d <= 8'hC0; 15'h05D9: d <= 8'hC0; 15'h05DA: d <= 8'hC0; 15'h05DB: d <= 8'hC0;
                15'h05DC: d <= 8'hC0; 15'h05DD: d <= 8'hC0; 15'h05DE: d <= 8'hC0; 15'h05DF: d <= 8'hC0;
                15'h05E0: d <= 8'hC0; 15'h05E1: d <= 8'hC0; 15'h05E2: d <= 8'hC0; 15'h05E3: d <= 8'hC0;
                15'h05E4: d <= 8'hC0; 15'h05E5: d <= 8'hC0; 15'h05E6: d <= 8'hC0; 15'h05E7: d <= 8'hC0;
                15'h05E8: d <= 8'hC0; 15'h05E9: d <= 8'hC0; 15'h05EA: d <= 8'hC0; 15'h05EB: d <= 8'hC0;
                15'h05EC: d <= 8'hC0; 15'h05ED: d <= 8'hC0; 15'h05EE: d <= 8'hC0; 15'h05EF: d <= 8'hC0;
                15'h05F0: d <= 8'hC0; 15'h05F1: d <= 8'hC0; 15'h05F2: d <= 8'hC0; 15'h05F3: d <= 8'hC0;
                15'h05F4: d <= 8'hC0; 15'h05F5: d <= 8'hC0; 15'h05F6: d <= 8'hC0; 15'h05F7: d <= 8'hC0;
                15'h05F8: d <= 8'hC0; 15'h05F9: d <= 8'hC0; 15'h05FA: d <= 8'hC0; 15'h05FB: d <= 8'hC0;
                15'h05FC: d <= 8'hC0; 15'h05FD: d <= 8'hC0; 15'h05FE: d <= 8'hC0; 15'h05FF: d <= 8'hC0;
                15'h0600: d <= 8'hC0; 15'h0601: d <= 8'hC0; 15'h0602: d <= 8'hC0; 15'h0603: d <= 8'hC0;
                15'h0604: d <= 8'hC0; 15'h0605: d <= 8'hC0; 15'h0606: d <= 8'hC0; 15'h0607: d <= 8'hC0;
                15'h0608: d <= 8'hC0; 15'h0609: d <= 8'hC0; 15'h060A: d <= 8'hC0; 15'h060B: d <= 8'hC0;
                15'h060C: d <= 8'hC0; 15'h060D: d <= 8'hC0; 15'h060E: d <= 8'hC0; 15'h060F: d <= 8'hC0;
                15'h0610: d <= 8'hC0; 15'h0611: d <= 8'hC0; 15'h0612: d <= 8'hC0; 15'h0613: d <= 8'hC0;
                15'h0614: d <= 8'hC0; 15'h0615: d <= 8'hC0; 15'h0616: d <= 8'hC0; 15'h0617: d <= 8'hC0;
                15'h0618: d <= 8'hC0; 15'h0619: d <= 8'hC0; 15'h061A: d <= 8'hC0; 15'h061B: d <= 8'hC0;
                15'h061C: d <= 8'hC0; 15'h061D: d <= 8'hC0; 15'h061E: d <= 8'hC0; 15'h061F: d <= 8'hC0;
                15'h0620: d <= 8'hC0; 15'h0621: d <= 8'hC0; 15'h0622: d <= 8'hC0; 15'h0623: d <= 8'hC0;
                15'h0624: d <= 8'hC0; 15'h0625: d <= 8'hC0; 15'h0626: d <= 8'hC0; 15'h0627: d <= 8'hC0;
                15'h0628: d <= 8'hC0; 15'h0629: d <= 8'hC0; 15'h062A: d <= 8'hC0; 15'h062B: d <= 8'hC0;
                15'h062C: d <= 8'hC0; 15'h062D: d <= 8'hC0; 15'h062E: d <= 8'hC0; 15'h062F: d <= 8'hC0;
                15'h0630: d <= 8'hC0; 15'h0631: d <= 8'hC0; 15'h0632: d <= 8'hC0; 15'h0633: d <= 8'hC0;
                15'h0634: d <= 8'hC0; 15'h0635: d <= 8'hC0; 15'h0636: d <= 8'hC0; 15'h0637: d <= 8'hC0;
                15'h0638: d <= 8'hC0; 15'h0639: d <= 8'hC0; 15'h063A: d <= 8'hC0; 15'h063B: d <= 8'hC0;
                15'h063C: d <= 8'hC0; 15'h063D: d <= 8'hC0; 15'h063E: d <= 8'hC0; 15'h063F: d <= 8'hC0;
                15'h0640: d <= 8'hC0; 15'h0641: d <= 8'hC0; 15'h0642: d <= 8'hC0; 15'h0643: d <= 8'hC0;
                15'h0644: d <= 8'hC0; 15'h0645: d <= 8'hC0; 15'h0646: d <= 8'hC0; 15'h0647: d <= 8'hC0;
                15'h0648: d <= 8'hC0; 15'h0649: d <= 8'hC0; 15'h064A: d <= 8'hC0; 15'h064B: d <= 8'hC0;
                15'h064C: d <= 8'hC0; 15'h064D: d <= 8'hC0; 15'h064E: d <= 8'hC0; 15'h064F: d <= 8'hC0;
                15'h0650: d <= 8'hC0; 15'h0651: d <= 8'hC0; 15'h0652: d <= 8'hC0; 15'h0653: d <= 8'hC0;
                15'h0654: d <= 8'hC0; 15'h0655: d <= 8'hC0; 15'h0656: d <= 8'hC0; 15'h0657: d <= 8'hC0;
                15'h0658: d <= 8'hC0; 15'h0659: d <= 8'hC0; 15'h065A: d <= 8'hC0; 15'h065B: d <= 8'hC0;
                15'h065C: d <= 8'hC0; 15'h065D: d <= 8'hC0; 15'h065E: d <= 8'hC0; 15'h065F: d <= 8'hC0;
                15'h0660: d <= 8'hC0; 15'h0661: d <= 8'hC0; 15'h0662: d <= 8'hC0; 15'h0663: d <= 8'hC0;
                15'h0664: d <= 8'hC0; 15'h0665: d <= 8'hC0; 15'h0666: d <= 8'hC0; 15'h0667: d <= 8'hC0;
                15'h0668: d <= 8'hC0; 15'h0669: d <= 8'hC0; 15'h066A: d <= 8'hC0; 15'h066B: d <= 8'hC0;
                15'h066C: d <= 8'hC0; 15'h066D: d <= 8'hC0; 15'h066E: d <= 8'hC0; 15'h066F: d <= 8'hC0;
                15'h0670: d <= 8'hC0; 15'h0671: d <= 8'hC0; 15'h0672: d <= 8'hC0; 15'h0673: d <= 8'hC0;
                15'h0674: d <= 8'hC0; 15'h0675: d <= 8'hC0; 15'h0676: d <= 8'hC0; 15'h0677: d <= 8'hC0;
                15'h0678: d <= 8'hC0; 15'h0679: d <= 8'hC0; 15'h067A: d <= 8'hC0; 15'h067B: d <= 8'hC0;
                15'h067C: d <= 8'hC0; 15'h067D: d <= 8'hC0; 15'h067E: d <= 8'hC0; 15'h067F: d <= 8'hC0;
                15'h0680: d <= 8'hC0; 15'h0681: d <= 8'hC0; 15'h0682: d <= 8'hC0; 15'h0683: d <= 8'hC0;
                15'h0684: d <= 8'hC0; 15'h0685: d <= 8'hC0; 15'h0686: d <= 8'hC0; 15'h0687: d <= 8'hC0;
                15'h0688: d <= 8'hC0; 15'h0689: d <= 8'hC0; 15'h068A: d <= 8'hC0; 15'h068B: d <= 8'hC0;
                15'h068C: d <= 8'hC0; 15'h068D: d <= 8'hC0; 15'h068E: d <= 8'hC0; 15'h068F: d <= 8'hC0;
                15'h0690: d <= 8'hC0; 15'h0691: d <= 8'hC0; 15'h0692: d <= 8'hC0; 15'h0693: d <= 8'hC0;
                15'h0694: d <= 8'hC0; 15'h0695: d <= 8'hC0; 15'h0696: d <= 8'hC0; 15'h0697: d <= 8'hC0;
                15'h0698: d <= 8'hC0; 15'h0699: d <= 8'hC0; 15'h069A: d <= 8'hC0; 15'h069B: d <= 8'hC0;
                15'h069C: d <= 8'hC0; 15'h069D: d <= 8'hC0; 15'h069E: d <= 8'hC0; 15'h069F: d <= 8'hC0;
                15'h06A0: d <= 8'hC0; 15'h06A1: d <= 8'hC0; 15'h06A2: d <= 8'hC0; 15'h06A3: d <= 8'hC0;
                15'h06A4: d <= 8'hC0; 15'h06A5: d <= 8'hC0; 15'h06A6: d <= 8'hC0; 15'h06A7: d <= 8'hC0;
                15'h06A8: d <= 8'hC0; 15'h06A9: d <= 8'hC0; 15'h06AA: d <= 8'hC0; 15'h06AB: d <= 8'hC0;
                15'h06AC: d <= 8'hC0; 15'h06AD: d <= 8'hC0; 15'h06AE: d <= 8'hC0; 15'h06AF: d <= 8'hC0;
                15'h06B0: d <= 8'hC0; 15'h06B1: d <= 8'hC0; 15'h06B2: d <= 8'hC0; 15'h06B3: d <= 8'hC0;
                15'h06B4: d <= 8'hC0; 15'h06B5: d <= 8'hC0; 15'h06B6: d <= 8'hC0; 15'h06B7: d <= 8'hC0;
                15'h06B8: d <= 8'hC0; 15'h06B9: d <= 8'hC0; 15'h06BA: d <= 8'hC0; 15'h06BB: d <= 8'hC0;
                15'h06BC: d <= 8'hC0; 15'h06BD: d <= 8'hC0; 15'h06BE: d <= 8'hC0; 15'h06BF: d <= 8'hC0;
                15'h06C0: d <= 8'hC0; 15'h06C1: d <= 8'hC0; 15'h06C2: d <= 8'hC0; 15'h06C3: d <= 8'hC0;
                15'h06C4: d <= 8'hC0; 15'h06C5: d <= 8'hC0; 15'h06C6: d <= 8'hC0; 15'h06C7: d <= 8'hC0;
                15'h06C8: d <= 8'hC0; 15'h06C9: d <= 8'hC0; 15'h06CA: d <= 8'hC0; 15'h06CB: d <= 8'hC0;
                15'h06CC: d <= 8'hC0; 15'h06CD: d <= 8'hC0; 15'h06CE: d <= 8'hC0; 15'h06CF: d <= 8'hC0;
                15'h06D0: d <= 8'hC0; 15'h06D1: d <= 8'hC0; 15'h06D2: d <= 8'hC0; 15'h06D3: d <= 8'hC0;
                15'h06D4: d <= 8'hC0; 15'h06D5: d <= 8'hC0; 15'h06D6: d <= 8'hC0; 15'h06D7: d <= 8'hC0;
                15'h06D8: d <= 8'hC0; 15'h06D9: d <= 8'hC0; 15'h06DA: d <= 8'hC0; 15'h06DB: d <= 8'hC0;
                15'h06DC: d <= 8'hC0; 15'h06DD: d <= 8'hC0; 15'h06DE: d <= 8'hC0; 15'h06DF: d <= 8'hC0;
                15'h06E0: d <= 8'hC0; 15'h06E1: d <= 8'hC0; 15'h06E2: d <= 8'hC0; 15'h06E3: d <= 8'hC0;
                15'h06E4: d <= 8'hC0; 15'h06E5: d <= 8'hC0; 15'h06E6: d <= 8'hC0; 15'h06E7: d <= 8'hC0;
                15'h06E8: d <= 8'hC0; 15'h06E9: d <= 8'hC0; 15'h06EA: d <= 8'hC0; 15'h06EB: d <= 8'hC0;
                15'h06EC: d <= 8'hC0; 15'h06ED: d <= 8'hC0; 15'h06EE: d <= 8'hC0; 15'h06EF: d <= 8'hC0;
                15'h06F0: d <= 8'hC0; 15'h06F1: d <= 8'hC0; 15'h06F2: d <= 8'hC0; 15'h06F3: d <= 8'hC0;
                15'h06F4: d <= 8'hC0; 15'h06F5: d <= 8'hC0; 15'h06F6: d <= 8'hC0; 15'h06F7: d <= 8'hC0;
                15'h06F8: d <= 8'hC0; 15'h06F9: d <= 8'hC0; 15'h06FA: d <= 8'hC0; 15'h06FB: d <= 8'hC0;
                15'h06FC: d <= 8'hC0; 15'h06FD: d <= 8'hC0; 15'h06FE: d <= 8'hC0; 15'h06FF: d <= 8'hC0;
                15'h0700: d <= 8'hC0; 15'h0701: d <= 8'hC0; 15'h0702: d <= 8'hC0; 15'h0703: d <= 8'hC0;
                15'h0704: d <= 8'hC0; 15'h0705: d <= 8'hC0; 15'h0706: d <= 8'hC0; 15'h0707: d <= 8'hC0;
                15'h0708: d <= 8'hC0; 15'h0709: d <= 8'hC0; 15'h070A: d <= 8'hC0; 15'h070B: d <= 8'hC0;
                15'h070C: d <= 8'hC0; 15'h070D: d <= 8'hC0; 15'h070E: d <= 8'hC0; 15'h070F: d <= 8'hC0;
                15'h0710: d <= 8'hC0; 15'h0711: d <= 8'hC0; 15'h0712: d <= 8'hC0; 15'h0713: d <= 8'hC0;
                15'h0714: d <= 8'hC0; 15'h0715: d <= 8'hC0; 15'h0716: d <= 8'hC0; 15'h0717: d <= 8'hC0;
                15'h0718: d <= 8'hC0; 15'h0719: d <= 8'hC0; 15'h071A: d <= 8'hC0; 15'h071B: d <= 8'hC0;
                15'h071C: d <= 8'hC0; 15'h071D: d <= 8'hC0; 15'h071E: d <= 8'hC0; 15'h071F: d <= 8'hC0;
                15'h0720: d <= 8'hC0; 15'h0721: d <= 8'hC0; 15'h0722: d <= 8'hC0; 15'h0723: d <= 8'hC0;
                15'h0724: d <= 8'hC0; 15'h0725: d <= 8'hC0; 15'h0726: d <= 8'hC0; 15'h0727: d <= 8'hC0;
                15'h0728: d <= 8'hC0; 15'h0729: d <= 8'hC0; 15'h072A: d <= 8'hC0; 15'h072B: d <= 8'hC0;
                15'h072C: d <= 8'hC0; 15'h072D: d <= 8'hC0; 15'h072E: d <= 8'hC0; 15'h072F: d <= 8'hC0;
                15'h0730: d <= 8'hC0; 15'h0731: d <= 8'hC0; 15'h0732: d <= 8'hC0; 15'h0733: d <= 8'hC0;
                15'h0734: d <= 8'hC0; 15'h0735: d <= 8'hC0; 15'h0736: d <= 8'hC0; 15'h0737: d <= 8'hC0;
                15'h0738: d <= 8'hC0; 15'h0739: d <= 8'hC0; 15'h073A: d <= 8'hC0; 15'h073B: d <= 8'hC0;
                15'h073C: d <= 8'hC0; 15'h073D: d <= 8'hC0; 15'h073E: d <= 8'hC0; 15'h073F: d <= 8'hC0;
                15'h0740: d <= 8'hC0; 15'h0741: d <= 8'hC0; 15'h0742: d <= 8'hC0; 15'h0743: d <= 8'hC0;
                15'h0744: d <= 8'hC0; 15'h0745: d <= 8'hC0; 15'h0746: d <= 8'hC0; 15'h0747: d <= 8'hC0;
                15'h0748: d <= 8'hC0; 15'h0749: d <= 8'hC0; 15'h074A: d <= 8'hC0; 15'h074B: d <= 8'hC0;
                15'h074C: d <= 8'hC0; 15'h074D: d <= 8'hC0; 15'h074E: d <= 8'hC0; 15'h074F: d <= 8'hC0;
                15'h0750: d <= 8'hC0; 15'h0751: d <= 8'hC0; 15'h0752: d <= 8'hC0; 15'h0753: d <= 8'hC0;
                15'h0754: d <= 8'hC0; 15'h0755: d <= 8'hC0; 15'h0756: d <= 8'hC0; 15'h0757: d <= 8'hC0;
                15'h0758: d <= 8'hC0; 15'h0759: d <= 8'hC0; 15'h075A: d <= 8'hC0; 15'h075B: d <= 8'hC0;
                15'h075C: d <= 8'hC0; 15'h075D: d <= 8'hC0; 15'h075E: d <= 8'hC0; 15'h075F: d <= 8'hC0;
                15'h0760: d <= 8'hC0; 15'h0761: d <= 8'hC0; 15'h0762: d <= 8'hC0; 15'h0763: d <= 8'hC0;
                15'h0764: d <= 8'hC0; 15'h0765: d <= 8'hC0; 15'h0766: d <= 8'hC0; 15'h0767: d <= 8'hC0;
                15'h0768: d <= 8'hC0; 15'h0769: d <= 8'hC0; 15'h076A: d <= 8'hC0; 15'h076B: d <= 8'hC0;
                15'h076C: d <= 8'hC0; 15'h076D: d <= 8'hC0; 15'h076E: d <= 8'hC0; 15'h076F: d <= 8'hC0;
                15'h0770: d <= 8'hC0; 15'h0771: d <= 8'hC0; 15'h0772: d <= 8'hC0; 15'h0773: d <= 8'hC0;
                15'h0774: d <= 8'hC0; 15'h0775: d <= 8'hC0; 15'h0776: d <= 8'hC0; 15'h0777: d <= 8'hC0;
                15'h0778: d <= 8'hC0; 15'h0779: d <= 8'hC0; 15'h077A: d <= 8'hC0; 15'h077B: d <= 8'hC0;
                15'h077C: d <= 8'hC0; 15'h077D: d <= 8'hC0; 15'h077E: d <= 8'hC0; 15'h077F: d <= 8'hC0;
                15'h0780: d <= 8'hC0; 15'h0781: d <= 8'hC0; 15'h0782: d <= 8'hC0; 15'h0783: d <= 8'hC0;
                15'h0784: d <= 8'hC0; 15'h0785: d <= 8'hC0; 15'h0786: d <= 8'hC0; 15'h0787: d <= 8'hC0;
                15'h0788: d <= 8'hC0; 15'h0789: d <= 8'hC0; 15'h078A: d <= 8'hC0; 15'h078B: d <= 8'hC0;
                15'h078C: d <= 8'hC0; 15'h078D: d <= 8'hC0; 15'h078E: d <= 8'hC0; 15'h078F: d <= 8'hC0;
                15'h0790: d <= 8'hC0; 15'h0791: d <= 8'hC0; 15'h0792: d <= 8'hC0; 15'h0793: d <= 8'hC0;
                15'h0794: d <= 8'hC0; 15'h0795: d <= 8'hC0; 15'h0796: d <= 8'hC0; 15'h0797: d <= 8'hC0;
                15'h0798: d <= 8'hC0; 15'h0799: d <= 8'hC0; 15'h079A: d <= 8'hC0; 15'h079B: d <= 8'hC0;
                15'h079C: d <= 8'hC0; 15'h079D: d <= 8'hC0; 15'h079E: d <= 8'hC0; 15'h079F: d <= 8'hC0;
                15'h07A0: d <= 8'hC0; 15'h07A1: d <= 8'hC0; 15'h07A2: d <= 8'hC0; 15'h07A3: d <= 8'hC0;
                15'h07A4: d <= 8'hC0; 15'h07A5: d <= 8'hC0; 15'h07A6: d <= 8'hC0; 15'h07A7: d <= 8'hC0;
                15'h07A8: d <= 8'hC0; 15'h07A9: d <= 8'hC0; 15'h07AA: d <= 8'hC0; 15'h07AB: d <= 8'hC0;
                15'h07AC: d <= 8'hC0; 15'h07AD: d <= 8'hC0; 15'h07AE: d <= 8'hC0; 15'h07AF: d <= 8'hC0;
                15'h07B0: d <= 8'hC0; 15'h07B1: d <= 8'hC0; 15'h07B2: d <= 8'hC0; 15'h07B3: d <= 8'hC0;
                15'h07B4: d <= 8'hC0; 15'h07B5: d <= 8'hC0; 15'h07B6: d <= 8'hC0; 15'h07B7: d <= 8'hC0;
                15'h07B8: d <= 8'hC0; 15'h07B9: d <= 8'hC0; 15'h07BA: d <= 8'hC0; 15'h07BB: d <= 8'hC0;
                15'h07BC: d <= 8'hC0; 15'h07BD: d <= 8'hC0; 15'h07BE: d <= 8'hC0; 15'h07BF: d <= 8'hC0;
                15'h07C0: d <= 8'hC0; 15'h07C1: d <= 8'hC0; 15'h07C2: d <= 8'hC0; 15'h07C3: d <= 8'hC0;
                15'h07C4: d <= 8'hC0; 15'h07C5: d <= 8'hC0; 15'h07C6: d <= 8'hC0; 15'h07C7: d <= 8'hC0;
                15'h07C8: d <= 8'hC0; 15'h07C9: d <= 8'hC0; 15'h07CA: d <= 8'hC0; 15'h07CB: d <= 8'hC0;
                15'h07CC: d <= 8'hC0; 15'h07CD: d <= 8'hC0; 15'h07CE: d <= 8'hC0; 15'h07CF: d <= 8'hC0;
                15'h07D0: d <= 8'hC0; 15'h07D1: d <= 8'hC0; 15'h07D2: d <= 8'hC0; 15'h07D3: d <= 8'hC0;
                15'h07D4: d <= 8'hC0; 15'h07D5: d <= 8'hC0; 15'h07D6: d <= 8'hC0; 15'h07D7: d <= 8'hC0;
                15'h07D8: d <= 8'hC0; 15'h07D9: d <= 8'hC0; 15'h07DA: d <= 8'hC0; 15'h07DB: d <= 8'hC0;
                15'h07DC: d <= 8'hC0; 15'h07DD: d <= 8'hC0; 15'h07DE: d <= 8'hC0; 15'h07DF: d <= 8'hC0;
                15'h07E0: d <= 8'hC0; 15'h07E1: d <= 8'hC0; 15'h07E2: d <= 8'hC0; 15'h07E3: d <= 8'hC0;
                15'h07E4: d <= 8'hC0; 15'h07E5: d <= 8'hC0; 15'h07E6: d <= 8'hC0; 15'h07E7: d <= 8'hC0;
                15'h07E8: d <= 8'hC0; 15'h07E9: d <= 8'hC0; 15'h07EA: d <= 8'hC0; 15'h07EB: d <= 8'hC0;
                15'h07EC: d <= 8'hC0; 15'h07ED: d <= 8'hC0; 15'h07EE: d <= 8'hC0; 15'h07EF: d <= 8'hC0;
                15'h07F0: d <= 8'hC0; 15'h07F1: d <= 8'hC0; 15'h07F2: d <= 8'hC0; 15'h07F3: d <= 8'hC0;
                15'h07F4: d <= 8'hC0; 15'h07F5: d <= 8'hC0; 15'h07F6: d <= 8'hC0; 15'h07F7: d <= 8'hC0;
                15'h07F8: d <= 8'hC0; 15'h07F9: d <= 8'hC0; 15'h07FA: d <= 8'hC0; 15'h07FB: d <= 8'hC0;
                15'h07FC: d <= 8'hC0; 15'h07FD: d <= 8'hC0; 15'h07FE: d <= 8'hC0; 15'h07FF: d <= 8'hC0;
                15'h0800: d <= 8'hC0; 15'h0801: d <= 8'hC0; 15'h0802: d <= 8'hC0; 15'h0803: d <= 8'hC0;
                15'h0804: d <= 8'hC0; 15'h0805: d <= 8'hC0; 15'h0806: d <= 8'hC0; 15'h0807: d <= 8'hC0;
                15'h0808: d <= 8'hC0; 15'h0809: d <= 8'hC0; 15'h080A: d <= 8'hC0; 15'h080B: d <= 8'hC0;
                15'h080C: d <= 8'hC0; 15'h080D: d <= 8'hC0; 15'h080E: d <= 8'hC0; 15'h080F: d <= 8'hC0;
                15'h0810: d <= 8'hC0; 15'h0811: d <= 8'hC0; 15'h0812: d <= 8'hC0; 15'h0813: d <= 8'hC0;
                15'h0814: d <= 8'hC0; 15'h0815: d <= 8'hC0; 15'h0816: d <= 8'hC0; 15'h0817: d <= 8'hC0;
                15'h0818: d <= 8'hC0; 15'h0819: d <= 8'hC0; 15'h081A: d <= 8'hC0; 15'h081B: d <= 8'hC0;
                15'h081C: d <= 8'hC0; 15'h081D: d <= 8'hC0; 15'h081E: d <= 8'hC0; 15'h081F: d <= 8'hC0;
                15'h0820: d <= 8'hC0; 15'h0821: d <= 8'hC0; 15'h0822: d <= 8'hC0; 15'h0823: d <= 8'hC0;
                15'h0824: d <= 8'hC0; 15'h0825: d <= 8'hC0; 15'h0826: d <= 8'hC0; 15'h0827: d <= 8'hC0;
                15'h0828: d <= 8'hC0; 15'h0829: d <= 8'hC0; 15'h082A: d <= 8'hC0; 15'h082B: d <= 8'hC0;
                15'h082C: d <= 8'hC0; 15'h082D: d <= 8'hC0; 15'h082E: d <= 8'hC0; 15'h082F: d <= 8'hC0;
                15'h0830: d <= 8'hC0; 15'h0831: d <= 8'hC0; 15'h0832: d <= 8'hC0; 15'h0833: d <= 8'hC0;
                15'h0834: d <= 8'hC0; 15'h0835: d <= 8'hC0; 15'h0836: d <= 8'hC0; 15'h0837: d <= 8'hC0;
                15'h0838: d <= 8'hC0; 15'h0839: d <= 8'hC0; 15'h083A: d <= 8'hC0; 15'h083B: d <= 8'hC0;
                15'h083C: d <= 8'hC0; 15'h083D: d <= 8'hC0; 15'h083E: d <= 8'hC0; 15'h083F: d <= 8'hC0;
                15'h0840: d <= 8'hC0; 15'h0841: d <= 8'hC0; 15'h0842: d <= 8'hC0; 15'h0843: d <= 8'hC0;
                15'h0844: d <= 8'hC0; 15'h0845: d <= 8'hC0; 15'h0846: d <= 8'hC0; 15'h0847: d <= 8'hC0;
                15'h0848: d <= 8'hC0; 15'h0849: d <= 8'hC0; 15'h084A: d <= 8'hC0; 15'h084B: d <= 8'hC0;
                15'h084C: d <= 8'hC0; 15'h084D: d <= 8'hC0; 15'h084E: d <= 8'hC0; 15'h084F: d <= 8'hC0;
                15'h0850: d <= 8'hC0; 15'h0851: d <= 8'hC0; 15'h0852: d <= 8'hC0; 15'h0853: d <= 8'hC0;
                15'h0854: d <= 8'hC0; 15'h0855: d <= 8'hC0; 15'h0856: d <= 8'hC0; 15'h0857: d <= 8'hC0;
                15'h0858: d <= 8'hC0; 15'h0859: d <= 8'hC0; 15'h085A: d <= 8'hC0; 15'h085B: d <= 8'hC0;
                15'h085C: d <= 8'hC0; 15'h085D: d <= 8'hC0; 15'h085E: d <= 8'hC0; 15'h085F: d <= 8'hC0;
                15'h0860: d <= 8'hC0; 15'h0861: d <= 8'hC0; 15'h0862: d <= 8'hC0; 15'h0863: d <= 8'hC0;
                15'h0864: d <= 8'hC0; 15'h0865: d <= 8'hC0; 15'h0866: d <= 8'hC0; 15'h0867: d <= 8'hC0;
                15'h0868: d <= 8'hC0; 15'h0869: d <= 8'hC0; 15'h086A: d <= 8'hC0; 15'h086B: d <= 8'hC0;
                15'h086C: d <= 8'hC0; 15'h086D: d <= 8'hC0; 15'h086E: d <= 8'hC0; 15'h086F: d <= 8'hC0;
                15'h0870: d <= 8'hC0; 15'h0871: d <= 8'hC0; 15'h0872: d <= 8'hC0; 15'h0873: d <= 8'hC0;
                15'h0874: d <= 8'hC0; 15'h0875: d <= 8'hC0; 15'h0876: d <= 8'hC0; 15'h0877: d <= 8'hC0;
                15'h0878: d <= 8'hC0; 15'h0879: d <= 8'hC0; 15'h087A: d <= 8'hC0; 15'h087B: d <= 8'hC0;
                15'h087C: d <= 8'hC0; 15'h087D: d <= 8'hC0; 15'h087E: d <= 8'hC0; 15'h087F: d <= 8'hC0;
                15'h0880: d <= 8'hC0; 15'h0881: d <= 8'hC0; 15'h0882: d <= 8'hC0; 15'h0883: d <= 8'hC0;
                15'h0884: d <= 8'hC0; 15'h0885: d <= 8'hC0; 15'h0886: d <= 8'hC0; 15'h0887: d <= 8'hC0;
                15'h0888: d <= 8'hC0; 15'h0889: d <= 8'hC0; 15'h088A: d <= 8'hC0; 15'h088B: d <= 8'hC0;
                15'h088C: d <= 8'hC0; 15'h088D: d <= 8'hC0; 15'h088E: d <= 8'hC0; 15'h088F: d <= 8'hC0;
                15'h0890: d <= 8'hC0; 15'h0891: d <= 8'hC0; 15'h0892: d <= 8'hC0; 15'h0893: d <= 8'hC0;
                15'h0894: d <= 8'hC0; 15'h0895: d <= 8'hC0; 15'h0896: d <= 8'hC0; 15'h0897: d <= 8'hC0;
                15'h0898: d <= 8'hC0; 15'h0899: d <= 8'hC0; 15'h089A: d <= 8'hC0; 15'h089B: d <= 8'hC0;
                15'h089C: d <= 8'hC0; 15'h089D: d <= 8'hC0; 15'h089E: d <= 8'hC0; 15'h089F: d <= 8'hC0;
                15'h08A0: d <= 8'hC0; 15'h08A1: d <= 8'hC0; 15'h08A2: d <= 8'hC0; 15'h08A3: d <= 8'hC0;
                15'h08A4: d <= 8'hC0; 15'h08A5: d <= 8'hC0; 15'h08A6: d <= 8'hC0; 15'h08A7: d <= 8'hC0;
                15'h08A8: d <= 8'hC0; 15'h08A9: d <= 8'hC0; 15'h08AA: d <= 8'hC0; 15'h08AB: d <= 8'hC0;
                15'h08AC: d <= 8'hC0; 15'h08AD: d <= 8'hC0; 15'h08AE: d <= 8'hC0; 15'h08AF: d <= 8'hC0;
                15'h08B0: d <= 8'hC0; 15'h08B1: d <= 8'hC0; 15'h08B2: d <= 8'hC0; 15'h08B3: d <= 8'hC0;
                15'h08B4: d <= 8'hC0; 15'h08B5: d <= 8'hC0; 15'h08B6: d <= 8'hC0; 15'h08B7: d <= 8'hC0;
                15'h08B8: d <= 8'hC0; 15'h08B9: d <= 8'hC0; 15'h08BA: d <= 8'hC0; 15'h08BB: d <= 8'hC0;
                15'h08BC: d <= 8'hC0; 15'h08BD: d <= 8'hC0; 15'h08BE: d <= 8'hC0; 15'h08BF: d <= 8'hC0;
                15'h08C0: d <= 8'hC0; 15'h08C1: d <= 8'hC0; 15'h08C2: d <= 8'hC0; 15'h08C3: d <= 8'hC0;
                15'h08C4: d <= 8'hC0; 15'h08C5: d <= 8'hC0; 15'h08C6: d <= 8'hC0; 15'h08C7: d <= 8'hC0;
                15'h08C8: d <= 8'hC0; 15'h08C9: d <= 8'hC0; 15'h08CA: d <= 8'hC0; 15'h08CB: d <= 8'hC0;
                15'h08CC: d <= 8'hC0; 15'h08CD: d <= 8'hC0; 15'h08CE: d <= 8'hC0; 15'h08CF: d <= 8'hC0;
                15'h08D0: d <= 8'hC0; 15'h08D1: d <= 8'hC0; 15'h08D2: d <= 8'hC0; 15'h08D3: d <= 8'hC0;
                15'h08D4: d <= 8'hC0; 15'h08D5: d <= 8'hC0; 15'h08D6: d <= 8'hC0; 15'h08D7: d <= 8'hC0;
                15'h08D8: d <= 8'hC0; 15'h08D9: d <= 8'hC0; 15'h08DA: d <= 8'hC0; 15'h08DB: d <= 8'hC0;
                15'h08DC: d <= 8'hC0; 15'h08DD: d <= 8'hC0; 15'h08DE: d <= 8'hC0; 15'h08DF: d <= 8'hC0;
                15'h08E0: d <= 8'hC0; 15'h08E1: d <= 8'hC0; 15'h08E2: d <= 8'hC0; 15'h08E3: d <= 8'hC0;
                15'h08E4: d <= 8'hC0; 15'h08E5: d <= 8'hC0; 15'h08E6: d <= 8'hC0; 15'h08E7: d <= 8'hC0;
                15'h08E8: d <= 8'hC0; 15'h08E9: d <= 8'hC0; 15'h08EA: d <= 8'hC0; 15'h08EB: d <= 8'hC0;
                15'h08EC: d <= 8'hC0; 15'h08ED: d <= 8'hC0; 15'h08EE: d <= 8'hC0; 15'h08EF: d <= 8'hC0;
                15'h08F0: d <= 8'hC0; 15'h08F1: d <= 8'hC0; 15'h08F2: d <= 8'hC0; 15'h08F3: d <= 8'hC0;
                15'h08F4: d <= 8'hC0; 15'h08F5: d <= 8'hC0; 15'h08F6: d <= 8'hC0; 15'h08F7: d <= 8'hC0;
                15'h08F8: d <= 8'hC0; 15'h08F9: d <= 8'hC0; 15'h08FA: d <= 8'hC0; 15'h08FB: d <= 8'hC0;
                15'h08FC: d <= 8'hC0; 15'h08FD: d <= 8'hC0; 15'h08FE: d <= 8'hC0; 15'h08FF: d <= 8'hC0;
                15'h0900: d <= 8'hC0; 15'h0901: d <= 8'hC0; 15'h0902: d <= 8'hC0; 15'h0903: d <= 8'hC0;
                15'h0904: d <= 8'hC0; 15'h0905: d <= 8'hC0; 15'h0906: d <= 8'hC0; 15'h0907: d <= 8'hC0;
                15'h0908: d <= 8'hC0; 15'h0909: d <= 8'hC0; 15'h090A: d <= 8'hC0; 15'h090B: d <= 8'hC0;
                15'h090C: d <= 8'hC0; 15'h090D: d <= 8'hC0; 15'h090E: d <= 8'hC0; 15'h090F: d <= 8'hC0;
                15'h0910: d <= 8'hC0; 15'h0911: d <= 8'hC0; 15'h0912: d <= 8'hC0; 15'h0913: d <= 8'hC0;
                15'h0914: d <= 8'hC0; 15'h0915: d <= 8'hC0; 15'h0916: d <= 8'hC0; 15'h0917: d <= 8'hC0;
                15'h0918: d <= 8'hC0; 15'h0919: d <= 8'hC0; 15'h091A: d <= 8'hC0; 15'h091B: d <= 8'hC0;
                15'h091C: d <= 8'hC0; 15'h091D: d <= 8'hC0; 15'h091E: d <= 8'hC0; 15'h091F: d <= 8'hC0;
                15'h0920: d <= 8'hC0; 15'h0921: d <= 8'hC0; 15'h0922: d <= 8'hC0; 15'h0923: d <= 8'hC0;
                15'h0924: d <= 8'hC0; 15'h0925: d <= 8'hC0; 15'h0926: d <= 8'hC0; 15'h0927: d <= 8'hC0;
                15'h0928: d <= 8'hC0; 15'h0929: d <= 8'hC0; 15'h092A: d <= 8'hC0; 15'h092B: d <= 8'hC0;
                15'h092C: d <= 8'hC0; 15'h092D: d <= 8'hC0; 15'h092E: d <= 8'hC0; 15'h092F: d <= 8'hC0;
                15'h0930: d <= 8'hC0; 15'h0931: d <= 8'hC0; 15'h0932: d <= 8'hC0; 15'h0933: d <= 8'hC0;
                15'h0934: d <= 8'hC0; 15'h0935: d <= 8'hC0; 15'h0936: d <= 8'hC0; 15'h0937: d <= 8'hC0;
                15'h0938: d <= 8'hC0; 15'h0939: d <= 8'hC0; 15'h093A: d <= 8'hC0; 15'h093B: d <= 8'hC0;
                15'h093C: d <= 8'hC0; 15'h093D: d <= 8'hC0; 15'h093E: d <= 8'hC0; 15'h093F: d <= 8'hC0;
                15'h0940: d <= 8'hC0; 15'h0941: d <= 8'hC0; 15'h0942: d <= 8'hC0; 15'h0943: d <= 8'hC0;
                15'h0944: d <= 8'hC0; 15'h0945: d <= 8'hC0; 15'h0946: d <= 8'hC0; 15'h0947: d <= 8'hC0;
                15'h0948: d <= 8'hC0; 15'h0949: d <= 8'hC0; 15'h094A: d <= 8'hC0; 15'h094B: d <= 8'hC0;
                15'h094C: d <= 8'hC0; 15'h094D: d <= 8'hC0; 15'h094E: d <= 8'hC0; 15'h094F: d <= 8'hC0;
                15'h0950: d <= 8'hC0; 15'h0951: d <= 8'hC0; 15'h0952: d <= 8'hC0; 15'h0953: d <= 8'hC0;
                15'h0954: d <= 8'hC0; 15'h0955: d <= 8'hC0; 15'h0956: d <= 8'hC0; 15'h0957: d <= 8'hC0;
                15'h0958: d <= 8'hC0; 15'h0959: d <= 8'hC0; 15'h095A: d <= 8'hC0; 15'h095B: d <= 8'hC0;
                15'h095C: d <= 8'hC0; 15'h095D: d <= 8'hC0; 15'h095E: d <= 8'hC0; 15'h095F: d <= 8'hC0;
                15'h0960: d <= 8'hC0; 15'h0961: d <= 8'hC0; 15'h0962: d <= 8'hC0; 15'h0963: d <= 8'hC0;
                15'h0964: d <= 8'hC0; 15'h0965: d <= 8'hC0; 15'h0966: d <= 8'hC0; 15'h0967: d <= 8'hC0;
                15'h0968: d <= 8'hC0; 15'h0969: d <= 8'hC0; 15'h096A: d <= 8'hC0; 15'h096B: d <= 8'hC0;
                15'h096C: d <= 8'hC0; 15'h096D: d <= 8'hC0; 15'h096E: d <= 8'hC0; 15'h096F: d <= 8'hC0;
                15'h0970: d <= 8'hC0; 15'h0971: d <= 8'hC0; 15'h0972: d <= 8'hC0; 15'h0973: d <= 8'hC0;
                15'h0974: d <= 8'hC0; 15'h0975: d <= 8'hC0; 15'h0976: d <= 8'hC0; 15'h0977: d <= 8'hC0;
                15'h0978: d <= 8'hC0; 15'h0979: d <= 8'hC0; 15'h097A: d <= 8'hC0; 15'h097B: d <= 8'hC0;
                15'h097C: d <= 8'hC0; 15'h097D: d <= 8'hC0; 15'h097E: d <= 8'hC0; 15'h097F: d <= 8'hC0;
                15'h0980: d <= 8'hC0; 15'h0981: d <= 8'hC0; 15'h0982: d <= 8'hC0; 15'h0983: d <= 8'hC0;
                15'h0984: d <= 8'hC0; 15'h0985: d <= 8'hC0; 15'h0986: d <= 8'hC0; 15'h0987: d <= 8'hC0;
                15'h0988: d <= 8'hC0; 15'h0989: d <= 8'hC0; 15'h098A: d <= 8'hC0; 15'h098B: d <= 8'hC0;
                15'h098C: d <= 8'hC0; 15'h098D: d <= 8'hC0; 15'h098E: d <= 8'hC0; 15'h098F: d <= 8'hC0;
                15'h0990: d <= 8'hC0; 15'h0991: d <= 8'hC0; 15'h0992: d <= 8'hC0; 15'h0993: d <= 8'hC0;
                15'h0994: d <= 8'hC0; 15'h0995: d <= 8'hC0; 15'h0996: d <= 8'hC0; 15'h0997: d <= 8'hC0;
                15'h0998: d <= 8'hC0; 15'h0999: d <= 8'hC0; 15'h099A: d <= 8'hC0; 15'h099B: d <= 8'hC0;
                15'h099C: d <= 8'hC0; 15'h099D: d <= 8'hC0; 15'h099E: d <= 8'hC0; 15'h099F: d <= 8'hC0;
                15'h09A0: d <= 8'hC0; 15'h09A1: d <= 8'hC0; 15'h09A2: d <= 8'hC0; 15'h09A3: d <= 8'hC0;
                15'h09A4: d <= 8'hC0; 15'h09A5: d <= 8'hC0; 15'h09A6: d <= 8'hC0; 15'h09A7: d <= 8'hC0;
                15'h09A8: d <= 8'hC0; 15'h09A9: d <= 8'hC0; 15'h09AA: d <= 8'hC0; 15'h09AB: d <= 8'hC0;
                15'h09AC: d <= 8'hC0; 15'h09AD: d <= 8'hC0; 15'h09AE: d <= 8'hC0; 15'h09AF: d <= 8'hC0;
                15'h09B0: d <= 8'hC0; 15'h09B1: d <= 8'hC0; 15'h09B2: d <= 8'hC0; 15'h09B3: d <= 8'hC0;
                15'h09B4: d <= 8'hC0; 15'h09B5: d <= 8'hC0; 15'h09B6: d <= 8'hC0; 15'h09B7: d <= 8'hC0;
                15'h09B8: d <= 8'hC0; 15'h09B9: d <= 8'hC0; 15'h09BA: d <= 8'hC0; 15'h09BB: d <= 8'hC0;
                15'h09BC: d <= 8'hC0; 15'h09BD: d <= 8'hC0; 15'h09BE: d <= 8'hC0; 15'h09BF: d <= 8'hC0;
                15'h09C0: d <= 8'hC0; 15'h09C1: d <= 8'hC0; 15'h09C2: d <= 8'hC0; 15'h09C3: d <= 8'hC0;
                15'h09C4: d <= 8'hC0; 15'h09C5: d <= 8'hC0; 15'h09C6: d <= 8'hC0; 15'h09C7: d <= 8'hC0;
                15'h09C8: d <= 8'hC0; 15'h09C9: d <= 8'hC0; 15'h09CA: d <= 8'hC0; 15'h09CB: d <= 8'hC0;
                15'h09CC: d <= 8'hC0; 15'h09CD: d <= 8'hC0; 15'h09CE: d <= 8'hC0; 15'h09CF: d <= 8'hC0;
                15'h09D0: d <= 8'hC0; 15'h09D1: d <= 8'hC0; 15'h09D2: d <= 8'hC0; 15'h09D3: d <= 8'hC0;
                15'h09D4: d <= 8'hC0; 15'h09D5: d <= 8'hC0; 15'h09D6: d <= 8'hC0; 15'h09D7: d <= 8'hC0;
                15'h09D8: d <= 8'hC0; 15'h09D9: d <= 8'hC0; 15'h09DA: d <= 8'hC0; 15'h09DB: d <= 8'hC0;
                15'h09DC: d <= 8'hC0; 15'h09DD: d <= 8'hC0; 15'h09DE: d <= 8'hC0; 15'h09DF: d <= 8'hC0;
                15'h09E0: d <= 8'hC0; 15'h09E1: d <= 8'hC0; 15'h09E2: d <= 8'hC0; 15'h09E3: d <= 8'hC0;
                15'h09E4: d <= 8'hC0; 15'h09E5: d <= 8'hC0; 15'h09E6: d <= 8'hC0; 15'h09E7: d <= 8'hC0;
                15'h09E8: d <= 8'hC0; 15'h09E9: d <= 8'hC0; 15'h09EA: d <= 8'hC0; 15'h09EB: d <= 8'hC0;
                15'h09EC: d <= 8'hC0; 15'h09ED: d <= 8'hC0; 15'h09EE: d <= 8'hC0; 15'h09EF: d <= 8'hC0;
                15'h09F0: d <= 8'hC0; 15'h09F1: d <= 8'hC0; 15'h09F2: d <= 8'hC0; 15'h09F3: d <= 8'hC0;
                15'h09F4: d <= 8'hC0; 15'h09F5: d <= 8'hC0; 15'h09F6: d <= 8'hC0; 15'h09F7: d <= 8'hC0;
                15'h09F8: d <= 8'hC0; 15'h09F9: d <= 8'hC0; 15'h09FA: d <= 8'hC0; 15'h09FB: d <= 8'hC0;
                15'h09FC: d <= 8'hC0; 15'h09FD: d <= 8'hC0; 15'h09FE: d <= 8'hC0; 15'h09FF: d <= 8'hC0;
                15'h0A00: d <= 8'hC0; 15'h0A01: d <= 8'hC0; 15'h0A02: d <= 8'hC0; 15'h0A03: d <= 8'hC0;
                15'h0A04: d <= 8'hC0; 15'h0A05: d <= 8'hC0; 15'h0A06: d <= 8'hC0; 15'h0A07: d <= 8'hC0;
                15'h0A08: d <= 8'hC0; 15'h0A09: d <= 8'hC0; 15'h0A0A: d <= 8'hC0; 15'h0A0B: d <= 8'hC0;
                15'h0A0C: d <= 8'hC0; 15'h0A0D: d <= 8'hC0; 15'h0A0E: d <= 8'hC0; 15'h0A0F: d <= 8'hC0;
                15'h0A10: d <= 8'hC0; 15'h0A11: d <= 8'hC0; 15'h0A12: d <= 8'hC0; 15'h0A13: d <= 8'hC0;
                15'h0A14: d <= 8'hC0; 15'h0A15: d <= 8'hC0; 15'h0A16: d <= 8'hC0; 15'h0A17: d <= 8'hC0;
                15'h0A18: d <= 8'hC0; 15'h0A19: d <= 8'hC0; 15'h0A1A: d <= 8'hC0; 15'h0A1B: d <= 8'hC0;
                15'h0A1C: d <= 8'hC0; 15'h0A1D: d <= 8'hC0; 15'h0A1E: d <= 8'hC0; 15'h0A1F: d <= 8'hC0;
                15'h0A20: d <= 8'hC0; 15'h0A21: d <= 8'hC0; 15'h0A22: d <= 8'hC0; 15'h0A23: d <= 8'hC0;
                15'h0A24: d <= 8'hC0; 15'h0A25: d <= 8'hC0; 15'h0A26: d <= 8'hC0; 15'h0A27: d <= 8'hC0;
                15'h0A28: d <= 8'hC0; 15'h0A29: d <= 8'hC0; 15'h0A2A: d <= 8'hC0; 15'h0A2B: d <= 8'hC0;
                15'h0A2C: d <= 8'hC0; 15'h0A2D: d <= 8'hC0; 15'h0A2E: d <= 8'hC0; 15'h0A2F: d <= 8'hC0;
                15'h0A30: d <= 8'hC0; 15'h0A31: d <= 8'hC0; 15'h0A32: d <= 8'hC0; 15'h0A33: d <= 8'hC0;
                15'h0A34: d <= 8'hC0; 15'h0A35: d <= 8'hC0; 15'h0A36: d <= 8'hC0; 15'h0A37: d <= 8'hC0;
                15'h0A38: d <= 8'hC0; 15'h0A39: d <= 8'hC0; 15'h0A3A: d <= 8'hC0; 15'h0A3B: d <= 8'hC0;
                15'h0A3C: d <= 8'hC0; 15'h0A3D: d <= 8'hC0; 15'h0A3E: d <= 8'hC0; 15'h0A3F: d <= 8'hC0;
                15'h0A40: d <= 8'hC0; 15'h0A41: d <= 8'hC0; 15'h0A42: d <= 8'hC0; 15'h0A43: d <= 8'hC0;
                15'h0A44: d <= 8'hC0; 15'h0A45: d <= 8'hC0; 15'h0A46: d <= 8'hC0; 15'h0A47: d <= 8'hC0;
                15'h0A48: d <= 8'hC0; 15'h0A49: d <= 8'hC0; 15'h0A4A: d <= 8'hC0; 15'h0A4B: d <= 8'hC0;
                15'h0A4C: d <= 8'hC0; 15'h0A4D: d <= 8'hC0; 15'h0A4E: d <= 8'hC0; 15'h0A4F: d <= 8'hC0;
                15'h0A50: d <= 8'hC0; 15'h0A51: d <= 8'hC0; 15'h0A52: d <= 8'hC0; 15'h0A53: d <= 8'hC0;
                15'h0A54: d <= 8'hC0; 15'h0A55: d <= 8'hC0; 15'h0A56: d <= 8'hC0; 15'h0A57: d <= 8'hC0;
                15'h0A58: d <= 8'hC0; 15'h0A59: d <= 8'hC0; 15'h0A5A: d <= 8'hC0; 15'h0A5B: d <= 8'hC0;
                15'h0A5C: d <= 8'hC0; 15'h0A5D: d <= 8'hC0; 15'h0A5E: d <= 8'hC0; 15'h0A5F: d <= 8'hC0;
                15'h0A60: d <= 8'hC0; 15'h0A61: d <= 8'hC0; 15'h0A62: d <= 8'hC0; 15'h0A63: d <= 8'hC0;
                15'h0A64: d <= 8'hC0; 15'h0A65: d <= 8'hC0; 15'h0A66: d <= 8'hC0; 15'h0A67: d <= 8'hC0;
                15'h0A68: d <= 8'hC0; 15'h0A69: d <= 8'hC0; 15'h0A6A: d <= 8'hC0; 15'h0A6B: d <= 8'hC0;
                15'h0A6C: d <= 8'hC0; 15'h0A6D: d <= 8'hC0; 15'h0A6E: d <= 8'hC0; 15'h0A6F: d <= 8'hC0;
                15'h0A70: d <= 8'hC0; 15'h0A71: d <= 8'hC0; 15'h0A72: d <= 8'hC0; 15'h0A73: d <= 8'hC0;
                15'h0A74: d <= 8'hC0; 15'h0A75: d <= 8'hC0; 15'h0A76: d <= 8'hC0; 15'h0A77: d <= 8'hC0;
                15'h0A78: d <= 8'hC0; 15'h0A79: d <= 8'hC0; 15'h0A7A: d <= 8'hC0; 15'h0A7B: d <= 8'hC0;
                15'h0A7C: d <= 8'hC0; 15'h0A7D: d <= 8'hC0; 15'h0A7E: d <= 8'hC0; 15'h0A7F: d <= 8'hC0;
                15'h0A80: d <= 8'hC0; 15'h0A81: d <= 8'hC0; 15'h0A82: d <= 8'hC0; 15'h0A83: d <= 8'hC0;
                15'h0A84: d <= 8'hC0; 15'h0A85: d <= 8'hC0; 15'h0A86: d <= 8'hC0; 15'h0A87: d <= 8'hC0;
                15'h0A88: d <= 8'hC0; 15'h0A89: d <= 8'hC0; 15'h0A8A: d <= 8'hC0; 15'h0A8B: d <= 8'hC0;
                15'h0A8C: d <= 8'hC0; 15'h0A8D: d <= 8'hC0; 15'h0A8E: d <= 8'hC0; 15'h0A8F: d <= 8'hC0;
                15'h0A90: d <= 8'hC0; 15'h0A91: d <= 8'hC0; 15'h0A92: d <= 8'hC0; 15'h0A93: d <= 8'hC0;
                15'h0A94: d <= 8'hC0; 15'h0A95: d <= 8'hC0; 15'h0A96: d <= 8'hC0; 15'h0A97: d <= 8'hC0;
                15'h0A98: d <= 8'hC0; 15'h0A99: d <= 8'hC0; 15'h0A9A: d <= 8'hC0; 15'h0A9B: d <= 8'hC0;
                15'h0A9C: d <= 8'hC0; 15'h0A9D: d <= 8'hC0; 15'h0A9E: d <= 8'hC0; 15'h0A9F: d <= 8'hC0;
                15'h0AA0: d <= 8'hC0; 15'h0AA1: d <= 8'hC0; 15'h0AA2: d <= 8'hC0; 15'h0AA3: d <= 8'hC0;
                15'h0AA4: d <= 8'hC0; 15'h0AA5: d <= 8'hC0; 15'h0AA6: d <= 8'hC0; 15'h0AA7: d <= 8'hC0;
                15'h0AA8: d <= 8'hC0; 15'h0AA9: d <= 8'hC0; 15'h0AAA: d <= 8'hC0; 15'h0AAB: d <= 8'hC0;
                15'h0AAC: d <= 8'hC0; 15'h0AAD: d <= 8'hC0; 15'h0AAE: d <= 8'hC0; 15'h0AAF: d <= 8'hC0;
                15'h0AB0: d <= 8'hC0; 15'h0AB1: d <= 8'hC0; 15'h0AB2: d <= 8'hC0; 15'h0AB3: d <= 8'hC0;
                15'h0AB4: d <= 8'hC0; 15'h0AB5: d <= 8'hC0; 15'h0AB6: d <= 8'hC0; 15'h0AB7: d <= 8'hC0;
                15'h0AB8: d <= 8'hC0; 15'h0AB9: d <= 8'hC0; 15'h0ABA: d <= 8'hC0; 15'h0ABB: d <= 8'hC0;
                15'h0ABC: d <= 8'hC0; 15'h0ABD: d <= 8'hC0; 15'h0ABE: d <= 8'hC0; 15'h0ABF: d <= 8'hC0;
                15'h0AC0: d <= 8'hC0; 15'h0AC1: d <= 8'hC0; 15'h0AC2: d <= 8'hC0; 15'h0AC3: d <= 8'hC0;
                15'h0AC4: d <= 8'hC0; 15'h0AC5: d <= 8'hC0; 15'h0AC6: d <= 8'hC0; 15'h0AC7: d <= 8'hC0;
                15'h0AC8: d <= 8'hC0; 15'h0AC9: d <= 8'hC0; 15'h0ACA: d <= 8'hC0; 15'h0ACB: d <= 8'hC0;
                15'h0ACC: d <= 8'hC0; 15'h0ACD: d <= 8'hC0; 15'h0ACE: d <= 8'hC0; 15'h0ACF: d <= 8'hC0;
                15'h0AD0: d <= 8'hC0; 15'h0AD1: d <= 8'hC0; 15'h0AD2: d <= 8'hC0; 15'h0AD3: d <= 8'hC0;
                15'h0AD4: d <= 8'hC0; 15'h0AD5: d <= 8'hC0; 15'h0AD6: d <= 8'hC0; 15'h0AD7: d <= 8'hC0;
                15'h0AD8: d <= 8'hC0; 15'h0AD9: d <= 8'hC0; 15'h0ADA: d <= 8'hC0; 15'h0ADB: d <= 8'hC0;
                15'h0ADC: d <= 8'hC0; 15'h0ADD: d <= 8'hC0; 15'h0ADE: d <= 8'hC0; 15'h0ADF: d <= 8'hC0;
                15'h0AE0: d <= 8'hC0; 15'h0AE1: d <= 8'hC0; 15'h0AE2: d <= 8'hC0; 15'h0AE3: d <= 8'hC0;
                15'h0AE4: d <= 8'hC0; 15'h0AE5: d <= 8'hC0; 15'h0AE6: d <= 8'hC0; 15'h0AE7: d <= 8'hC0;
                15'h0AE8: d <= 8'hC0; 15'h0AE9: d <= 8'hC0; 15'h0AEA: d <= 8'hC0; 15'h0AEB: d <= 8'hC0;
                15'h0AEC: d <= 8'hC0; 15'h0AED: d <= 8'hC0; 15'h0AEE: d <= 8'hC0; 15'h0AEF: d <= 8'hC0;
                15'h0AF0: d <= 8'hC0; 15'h0AF1: d <= 8'hC0; 15'h0AF2: d <= 8'hC0; 15'h0AF3: d <= 8'hC0;
                15'h0AF4: d <= 8'hC0; 15'h0AF5: d <= 8'hC0; 15'h0AF6: d <= 8'hC0; 15'h0AF7: d <= 8'hC0;
                15'h0AF8: d <= 8'hC0; 15'h0AF9: d <= 8'hC0; 15'h0AFA: d <= 8'hC0; 15'h0AFB: d <= 8'hC0;
                15'h0AFC: d <= 8'hC0; 15'h0AFD: d <= 8'hC0; 15'h0AFE: d <= 8'hC0; 15'h0AFF: d <= 8'hC0;
                15'h0B00: d <= 8'hC0; 15'h0B01: d <= 8'hC0; 15'h0B02: d <= 8'hC0; 15'h0B03: d <= 8'hC0;
                15'h0B04: d <= 8'hC0; 15'h0B05: d <= 8'hC0; 15'h0B06: d <= 8'hC0; 15'h0B07: d <= 8'hC0;
                15'h0B08: d <= 8'hC0; 15'h0B09: d <= 8'hC0; 15'h0B0A: d <= 8'hC0; 15'h0B0B: d <= 8'hC0;
                15'h0B0C: d <= 8'hC0; 15'h0B0D: d <= 8'hC0; 15'h0B0E: d <= 8'hC0; 15'h0B0F: d <= 8'hC0;
                15'h0B10: d <= 8'hC0; 15'h0B11: d <= 8'hC0; 15'h0B12: d <= 8'hC0; 15'h0B13: d <= 8'hC0;
                15'h0B14: d <= 8'hC0; 15'h0B15: d <= 8'hC0; 15'h0B16: d <= 8'hC0; 15'h0B17: d <= 8'hC0;
                15'h0B18: d <= 8'hC0; 15'h0B19: d <= 8'hC0; 15'h0B1A: d <= 8'hC0; 15'h0B1B: d <= 8'hC0;
                15'h0B1C: d <= 8'hC0; 15'h0B1D: d <= 8'hC0; 15'h0B1E: d <= 8'hC0; 15'h0B1F: d <= 8'hC0;
                15'h0B20: d <= 8'hC0; 15'h0B21: d <= 8'hC0; 15'h0B22: d <= 8'hC0; 15'h0B23: d <= 8'hC0;
                15'h0B24: d <= 8'hC0; 15'h0B25: d <= 8'hC0; 15'h0B26: d <= 8'hC0; 15'h0B27: d <= 8'hC0;
                15'h0B28: d <= 8'hC0; 15'h0B29: d <= 8'hC0; 15'h0B2A: d <= 8'hC0; 15'h0B2B: d <= 8'hC0;
                15'h0B2C: d <= 8'hC0; 15'h0B2D: d <= 8'hC0; 15'h0B2E: d <= 8'hC0; 15'h0B2F: d <= 8'hC0;
                15'h0B30: d <= 8'hC0; 15'h0B31: d <= 8'hC0; 15'h0B32: d <= 8'hC0; 15'h0B33: d <= 8'hC0;
                15'h0B34: d <= 8'hC0; 15'h0B35: d <= 8'hC0; 15'h0B36: d <= 8'hC0; 15'h0B37: d <= 8'hC0;
                15'h0B38: d <= 8'hC0; 15'h0B39: d <= 8'hC0; 15'h0B3A: d <= 8'hC0; 15'h0B3B: d <= 8'hC0;
                15'h0B3C: d <= 8'hC0; 15'h0B3D: d <= 8'hC0; 15'h0B3E: d <= 8'hC0; 15'h0B3F: d <= 8'hC0;
                15'h0B40: d <= 8'hC0; 15'h0B41: d <= 8'hC0; 15'h0B42: d <= 8'hC0; 15'h0B43: d <= 8'hC0;
                15'h0B44: d <= 8'hC0; 15'h0B45: d <= 8'hC0; 15'h0B46: d <= 8'hC0; 15'h0B47: d <= 8'hC0;
                15'h0B48: d <= 8'hC0; 15'h0B49: d <= 8'hC0; 15'h0B4A: d <= 8'hC0; 15'h0B4B: d <= 8'hC0;
                15'h0B4C: d <= 8'hC0; 15'h0B4D: d <= 8'hC0; 15'h0B4E: d <= 8'hC0; 15'h0B4F: d <= 8'hC0;
                15'h0B50: d <= 8'hC0; 15'h0B51: d <= 8'hC0; 15'h0B52: d <= 8'hC0; 15'h0B53: d <= 8'hC0;
                15'h0B54: d <= 8'hC0; 15'h0B55: d <= 8'hC0; 15'h0B56: d <= 8'hC0; 15'h0B57: d <= 8'hC0;
                15'h0B58: d <= 8'hC0; 15'h0B59: d <= 8'hC0; 15'h0B5A: d <= 8'hC0; 15'h0B5B: d <= 8'hC0;
                15'h0B5C: d <= 8'hC0; 15'h0B5D: d <= 8'hC0; 15'h0B5E: d <= 8'hC0; 15'h0B5F: d <= 8'hC0;
                15'h0B60: d <= 8'hC0; 15'h0B61: d <= 8'hC0; 15'h0B62: d <= 8'hC0; 15'h0B63: d <= 8'hC0;
                15'h0B64: d <= 8'hC0; 15'h0B65: d <= 8'hC0; 15'h0B66: d <= 8'hC0; 15'h0B67: d <= 8'hC0;
                15'h0B68: d <= 8'hC0; 15'h0B69: d <= 8'hC0; 15'h0B6A: d <= 8'hC0; 15'h0B6B: d <= 8'hC0;
                15'h0B6C: d <= 8'hC0; 15'h0B6D: d <= 8'hC0; 15'h0B6E: d <= 8'hC0; 15'h0B6F: d <= 8'hC0;
                15'h0B70: d <= 8'hC0; 15'h0B71: d <= 8'hC0; 15'h0B72: d <= 8'hC0; 15'h0B73: d <= 8'hC0;
                15'h0B74: d <= 8'hC0; 15'h0B75: d <= 8'hC0; 15'h0B76: d <= 8'hC0; 15'h0B77: d <= 8'hC0;
                15'h0B78: d <= 8'hC0; 15'h0B79: d <= 8'hC0; 15'h0B7A: d <= 8'hC0; 15'h0B7B: d <= 8'hC0;
                15'h0B7C: d <= 8'hC0; 15'h0B7D: d <= 8'hC0; 15'h0B7E: d <= 8'hC0; 15'h0B7F: d <= 8'hC0;
                15'h0B80: d <= 8'hC0; 15'h0B81: d <= 8'hC0; 15'h0B82: d <= 8'hC0; 15'h0B83: d <= 8'hC0;
                15'h0B84: d <= 8'hC0; 15'h0B85: d <= 8'hC0; 15'h0B86: d <= 8'hC0; 15'h0B87: d <= 8'hC0;
                15'h0B88: d <= 8'hC0; 15'h0B89: d <= 8'hC0; 15'h0B8A: d <= 8'hC0; 15'h0B8B: d <= 8'hC0;
                15'h0B8C: d <= 8'hC0; 15'h0B8D: d <= 8'hC0; 15'h0B8E: d <= 8'hC0; 15'h0B8F: d <= 8'hC0;
                15'h0B90: d <= 8'hC0; 15'h0B91: d <= 8'hC0; 15'h0B92: d <= 8'hC0; 15'h0B93: d <= 8'hC0;
                15'h0B94: d <= 8'hC0; 15'h0B95: d <= 8'hC0; 15'h0B96: d <= 8'hC0; 15'h0B97: d <= 8'hC0;
                15'h0B98: d <= 8'hC0; 15'h0B99: d <= 8'hC0; 15'h0B9A: d <= 8'hC0; 15'h0B9B: d <= 8'hC0;
                15'h0B9C: d <= 8'hC0; 15'h0B9D: d <= 8'hC0; 15'h0B9E: d <= 8'hC0; 15'h0B9F: d <= 8'hC0;
                15'h0BA0: d <= 8'hC0; 15'h0BA1: d <= 8'hC0; 15'h0BA2: d <= 8'hC0; 15'h0BA3: d <= 8'hC0;
                15'h0BA4: d <= 8'hC0; 15'h0BA5: d <= 8'hC0; 15'h0BA6: d <= 8'hC0; 15'h0BA7: d <= 8'hC0;
                15'h0BA8: d <= 8'hC0; 15'h0BA9: d <= 8'hC0; 15'h0BAA: d <= 8'hC0; 15'h0BAB: d <= 8'hC0;
                15'h0BAC: d <= 8'hC0; 15'h0BAD: d <= 8'hC0; 15'h0BAE: d <= 8'hC0; 15'h0BAF: d <= 8'hC0;
                15'h0BB0: d <= 8'hC0; 15'h0BB1: d <= 8'hC0; 15'h0BB2: d <= 8'hC0; 15'h0BB3: d <= 8'hC0;
                15'h0BB4: d <= 8'hC0; 15'h0BB5: d <= 8'hC0; 15'h0BB6: d <= 8'hC0; 15'h0BB7: d <= 8'hC0;
                15'h0BB8: d <= 8'hC0; 15'h0BB9: d <= 8'hC0; 15'h0BBA: d <= 8'hC0; 15'h0BBB: d <= 8'hC0;
                15'h0BBC: d <= 8'hC0; 15'h0BBD: d <= 8'hC0; 15'h0BBE: d <= 8'hC0; 15'h0BBF: d <= 8'hC0;
                15'h0BC0: d <= 8'hC0; 15'h0BC1: d <= 8'hC0; 15'h0BC2: d <= 8'hC0; 15'h0BC3: d <= 8'hC0;
                15'h0BC4: d <= 8'hC0; 15'h0BC5: d <= 8'hC0; 15'h0BC6: d <= 8'hC0; 15'h0BC7: d <= 8'hC0;
                15'h0BC8: d <= 8'hC0; 15'h0BC9: d <= 8'hC0; 15'h0BCA: d <= 8'hC0; 15'h0BCB: d <= 8'hC0;
                15'h0BCC: d <= 8'hC0; 15'h0BCD: d <= 8'hC0; 15'h0BCE: d <= 8'hC0; 15'h0BCF: d <= 8'hC0;
                15'h0BD0: d <= 8'hC0; 15'h0BD1: d <= 8'hC0; 15'h0BD2: d <= 8'hC0; 15'h0BD3: d <= 8'hC0;
                15'h0BD4: d <= 8'hC0; 15'h0BD5: d <= 8'hC0; 15'h0BD6: d <= 8'hC0; 15'h0BD7: d <= 8'hC0;
                15'h0BD8: d <= 8'hC0; 15'h0BD9: d <= 8'hC0; 15'h0BDA: d <= 8'hC0; 15'h0BDB: d <= 8'hC0;
                15'h0BDC: d <= 8'hC0; 15'h0BDD: d <= 8'hC0; 15'h0BDE: d <= 8'hC0; 15'h0BDF: d <= 8'hC0;
                15'h0BE0: d <= 8'hC0; 15'h0BE1: d <= 8'hC0; 15'h0BE2: d <= 8'hC0; 15'h0BE3: d <= 8'hC0;
                15'h0BE4: d <= 8'hC0; 15'h0BE5: d <= 8'hC0; 15'h0BE6: d <= 8'hC0; 15'h0BE7: d <= 8'hC0;
                15'h0BE8: d <= 8'hC0; 15'h0BE9: d <= 8'hC0; 15'h0BEA: d <= 8'hC0; 15'h0BEB: d <= 8'hC0;
                15'h0BEC: d <= 8'hC0; 15'h0BED: d <= 8'hC0; 15'h0BEE: d <= 8'hC0; 15'h0BEF: d <= 8'hC0;
                15'h0BF0: d <= 8'hC0; 15'h0BF1: d <= 8'hC0; 15'h0BF2: d <= 8'hC0; 15'h0BF3: d <= 8'hC0;
                15'h0BF4: d <= 8'hC0; 15'h0BF5: d <= 8'hC0; 15'h0BF6: d <= 8'hC0; 15'h0BF7: d <= 8'hC0;
                15'h0BF8: d <= 8'hC0; 15'h0BF9: d <= 8'hC0; 15'h0BFA: d <= 8'hC0; 15'h0BFB: d <= 8'hC0;
                15'h0BFC: d <= 8'hC0; 15'h0BFD: d <= 8'hC0; 15'h0BFE: d <= 8'hC0; 15'h0BFF: d <= 8'hC0;
                15'h0C00: d <= 8'hC0; 15'h0C01: d <= 8'hC0; 15'h0C02: d <= 8'hC0; 15'h0C03: d <= 8'hC0;
                15'h0C04: d <= 8'hC0; 15'h0C05: d <= 8'hC0; 15'h0C06: d <= 8'hC0; 15'h0C07: d <= 8'hC0;
                15'h0C08: d <= 8'hC0; 15'h0C09: d <= 8'hC0; 15'h0C0A: d <= 8'hC0; 15'h0C0B: d <= 8'hC0;
                15'h0C0C: d <= 8'hC0; 15'h0C0D: d <= 8'hC0; 15'h0C0E: d <= 8'hC0; 15'h0C0F: d <= 8'hC0;
                15'h0C10: d <= 8'hC0; 15'h0C11: d <= 8'hC0; 15'h0C12: d <= 8'hC0; 15'h0C13: d <= 8'hC0;
                15'h0C14: d <= 8'hC0; 15'h0C15: d <= 8'hC0; 15'h0C16: d <= 8'hC0; 15'h0C17: d <= 8'hC0;
                15'h0C18: d <= 8'hC0; 15'h0C19: d <= 8'hC0; 15'h0C1A: d <= 8'hC0; 15'h0C1B: d <= 8'hC0;
                15'h0C1C: d <= 8'hC0; 15'h0C1D: d <= 8'hC0; 15'h0C1E: d <= 8'hC0; 15'h0C1F: d <= 8'hC0;
                15'h0C20: d <= 8'hC0; 15'h0C21: d <= 8'hC0; 15'h0C22: d <= 8'hC0; 15'h0C23: d <= 8'hC0;
                15'h0C24: d <= 8'hC0; 15'h0C25: d <= 8'hC0; 15'h0C26: d <= 8'hC0; 15'h0C27: d <= 8'hC0;
                15'h0C28: d <= 8'hC0; 15'h0C29: d <= 8'hC0; 15'h0C2A: d <= 8'hC0; 15'h0C2B: d <= 8'hC0;
                15'h0C2C: d <= 8'hC0; 15'h0C2D: d <= 8'hC0; 15'h0C2E: d <= 8'hC0; 15'h0C2F: d <= 8'hC0;
                15'h0C30: d <= 8'hC0; 15'h0C31: d <= 8'hC0; 15'h0C32: d <= 8'hC0; 15'h0C33: d <= 8'hC0;
                15'h0C34: d <= 8'hC0; 15'h0C35: d <= 8'hC0; 15'h0C36: d <= 8'hC0; 15'h0C37: d <= 8'hC0;
                15'h0C38: d <= 8'hC0; 15'h0C39: d <= 8'hC0; 15'h0C3A: d <= 8'hC0; 15'h0C3B: d <= 8'hC0;
                15'h0C3C: d <= 8'hC0; 15'h0C3D: d <= 8'hC0; 15'h0C3E: d <= 8'hC0; 15'h0C3F: d <= 8'hC0;
                15'h0C40: d <= 8'hC0; 15'h0C41: d <= 8'hC0; 15'h0C42: d <= 8'hC0; 15'h0C43: d <= 8'hC0;
                15'h0C44: d <= 8'hC0; 15'h0C45: d <= 8'hC0; 15'h0C46: d <= 8'hC0; 15'h0C47: d <= 8'hC0;
                15'h0C48: d <= 8'hC0; 15'h0C49: d <= 8'hC0; 15'h0C4A: d <= 8'hC0; 15'h0C4B: d <= 8'hC0;
                15'h0C4C: d <= 8'hC0; 15'h0C4D: d <= 8'hC0; 15'h0C4E: d <= 8'hC0; 15'h0C4F: d <= 8'hC0;
                15'h0C50: d <= 8'hC0; 15'h0C51: d <= 8'hC0; 15'h0C52: d <= 8'hC0; 15'h0C53: d <= 8'hC0;
                15'h0C54: d <= 8'hC0; 15'h0C55: d <= 8'hC0; 15'h0C56: d <= 8'hC0; 15'h0C57: d <= 8'hC0;
                15'h0C58: d <= 8'hC0; 15'h0C59: d <= 8'hC0; 15'h0C5A: d <= 8'hC0; 15'h0C5B: d <= 8'hC0;
                15'h0C5C: d <= 8'hC0; 15'h0C5D: d <= 8'hC0; 15'h0C5E: d <= 8'hC0; 15'h0C5F: d <= 8'hC0;
                15'h0C60: d <= 8'hC0; 15'h0C61: d <= 8'hC0; 15'h0C62: d <= 8'hC0; 15'h0C63: d <= 8'hC0;
                15'h0C64: d <= 8'hC0; 15'h0C65: d <= 8'hC0; 15'h0C66: d <= 8'hC0; 15'h0C67: d <= 8'hC0;
                15'h0C68: d <= 8'hC0; 15'h0C69: d <= 8'hC0; 15'h0C6A: d <= 8'hC0; 15'h0C6B: d <= 8'hC0;
                15'h0C6C: d <= 8'hC0; 15'h0C6D: d <= 8'hC0; 15'h0C6E: d <= 8'hC0; 15'h0C6F: d <= 8'hC0;
                15'h0C70: d <= 8'hC0; 15'h0C71: d <= 8'hC0; 15'h0C72: d <= 8'hC0; 15'h0C73: d <= 8'hC0;
                15'h0C74: d <= 8'hC0; 15'h0C75: d <= 8'hC0; 15'h0C76: d <= 8'hC0; 15'h0C77: d <= 8'hC0;
                15'h0C78: d <= 8'hC0; 15'h0C79: d <= 8'hC0; 15'h0C7A: d <= 8'hC0; 15'h0C7B: d <= 8'hC0;
                15'h0C7C: d <= 8'hC0; 15'h0C7D: d <= 8'hC0; 15'h0C7E: d <= 8'hC0; 15'h0C7F: d <= 8'hC0;
                15'h0C80: d <= 8'hC0; 15'h0C81: d <= 8'hC0; 15'h0C82: d <= 8'hC0; 15'h0C83: d <= 8'hC0;
                15'h0C84: d <= 8'hC0; 15'h0C85: d <= 8'hC0; 15'h0C86: d <= 8'hC0; 15'h0C87: d <= 8'hC0;
                15'h0C88: d <= 8'hC0; 15'h0C89: d <= 8'hC0; 15'h0C8A: d <= 8'hC0; 15'h0C8B: d <= 8'hC0;
                15'h0C8C: d <= 8'hC0; 15'h0C8D: d <= 8'hC0; 15'h0C8E: d <= 8'hC0; 15'h0C8F: d <= 8'hC0;
                15'h0C90: d <= 8'hC0; 15'h0C91: d <= 8'hC0; 15'h0C92: d <= 8'hC0; 15'h0C93: d <= 8'hC0;
                15'h0C94: d <= 8'hC0; 15'h0C95: d <= 8'hC0; 15'h0C96: d <= 8'hC0; 15'h0C97: d <= 8'hC0;
                15'h0C98: d <= 8'hC0; 15'h0C99: d <= 8'hC0; 15'h0C9A: d <= 8'hC0; 15'h0C9B: d <= 8'hC0;
                15'h0C9C: d <= 8'hC0; 15'h0C9D: d <= 8'hC0; 15'h0C9E: d <= 8'hC0; 15'h0C9F: d <= 8'hC0;
                15'h0CA0: d <= 8'hC0; 15'h0CA1: d <= 8'hC0; 15'h0CA2: d <= 8'hC0; 15'h0CA3: d <= 8'hC0;
                15'h0CA4: d <= 8'hC0; 15'h0CA5: d <= 8'hC0; 15'h0CA6: d <= 8'hC0; 15'h0CA7: d <= 8'hC0;
                15'h0CA8: d <= 8'hC0; 15'h0CA9: d <= 8'hC0; 15'h0CAA: d <= 8'hC0; 15'h0CAB: d <= 8'hC0;
                15'h0CAC: d <= 8'hC0; 15'h0CAD: d <= 8'hC0; 15'h0CAE: d <= 8'hC0; 15'h0CAF: d <= 8'hC0;
                15'h0CB0: d <= 8'hC0; 15'h0CB1: d <= 8'hC0; 15'h0CB2: d <= 8'hC0; 15'h0CB3: d <= 8'hC0;
                15'h0CB4: d <= 8'hC0; 15'h0CB5: d <= 8'hC0; 15'h0CB6: d <= 8'hC0; 15'h0CB7: d <= 8'hC0;
                15'h0CB8: d <= 8'hC0; 15'h0CB9: d <= 8'hC0; 15'h0CBA: d <= 8'hC0; 15'h0CBB: d <= 8'hC0;
                15'h0CBC: d <= 8'hC0; 15'h0CBD: d <= 8'hC0; 15'h0CBE: d <= 8'hC0; 15'h0CBF: d <= 8'hC0;
                15'h0CC0: d <= 8'hC0; 15'h0CC1: d <= 8'hC0; 15'h0CC2: d <= 8'hC0; 15'h0CC3: d <= 8'hC0;
                15'h0CC4: d <= 8'hC0; 15'h0CC5: d <= 8'hC0; 15'h0CC6: d <= 8'hC0; 15'h0CC7: d <= 8'hC0;
                15'h0CC8: d <= 8'hC0; 15'h0CC9: d <= 8'hC0; 15'h0CCA: d <= 8'hC0; 15'h0CCB: d <= 8'hC0;
                15'h0CCC: d <= 8'hC0; 15'h0CCD: d <= 8'hC0; 15'h0CCE: d <= 8'hC0; 15'h0CCF: d <= 8'hC0;
                15'h0CD0: d <= 8'hC0; 15'h0CD1: d <= 8'hC0; 15'h0CD2: d <= 8'hC0; 15'h0CD3: d <= 8'hC0;
                15'h0CD4: d <= 8'hC0; 15'h0CD5: d <= 8'hC0; 15'h0CD6: d <= 8'hC0; 15'h0CD7: d <= 8'hC0;
                15'h0CD8: d <= 8'hC0; 15'h0CD9: d <= 8'hC0; 15'h0CDA: d <= 8'hC0; 15'h0CDB: d <= 8'hC0;
                15'h0CDC: d <= 8'hC0; 15'h0CDD: d <= 8'hC0; 15'h0CDE: d <= 8'hC0; 15'h0CDF: d <= 8'hC0;
                15'h0CE0: d <= 8'hC0; 15'h0CE1: d <= 8'hC0; 15'h0CE2: d <= 8'hC0; 15'h0CE3: d <= 8'hC0;
                15'h0CE4: d <= 8'hC0; 15'h0CE5: d <= 8'hC0; 15'h0CE6: d <= 8'hC0; 15'h0CE7: d <= 8'hC0;
                15'h0CE8: d <= 8'hC0; 15'h0CE9: d <= 8'hC0; 15'h0CEA: d <= 8'hC0; 15'h0CEB: d <= 8'hC0;
                15'h0CEC: d <= 8'hC0; 15'h0CED: d <= 8'hC0; 15'h0CEE: d <= 8'hC0; 15'h0CEF: d <= 8'hC0;
                15'h0CF0: d <= 8'hC0; 15'h0CF1: d <= 8'hC0; 15'h0CF2: d <= 8'hC0; 15'h0CF3: d <= 8'hC0;
                15'h0CF4: d <= 8'hC0; 15'h0CF5: d <= 8'hC0; 15'h0CF6: d <= 8'hC0; 15'h0CF7: d <= 8'hC0;
                15'h0CF8: d <= 8'hC0; 15'h0CF9: d <= 8'hC0; 15'h0CFA: d <= 8'hC0; 15'h0CFB: d <= 8'hC0;
                15'h0CFC: d <= 8'hC0; 15'h0CFD: d <= 8'hC0; 15'h0CFE: d <= 8'hC0; 15'h0CFF: d <= 8'hC0;
                15'h0D00: d <= 8'hC0; 15'h0D01: d <= 8'hC0; 15'h0D02: d <= 8'hC0; 15'h0D03: d <= 8'hC0;
                15'h0D04: d <= 8'hC0; 15'h0D05: d <= 8'hC0; 15'h0D06: d <= 8'hC0; 15'h0D07: d <= 8'hC0;
                15'h0D08: d <= 8'hC0; 15'h0D09: d <= 8'hC0; 15'h0D0A: d <= 8'hC0; 15'h0D0B: d <= 8'hC0;
                15'h0D0C: d <= 8'hC0; 15'h0D0D: d <= 8'hC0; 15'h0D0E: d <= 8'hC0; 15'h0D0F: d <= 8'hC0;
                15'h0D10: d <= 8'hC0; 15'h0D11: d <= 8'hC0; 15'h0D12: d <= 8'hC0; 15'h0D13: d <= 8'hC0;
                15'h0D14: d <= 8'hC0; 15'h0D15: d <= 8'hC0; 15'h0D16: d <= 8'hC0; 15'h0D17: d <= 8'hC0;
                15'h0D18: d <= 8'hC0; 15'h0D19: d <= 8'hC0; 15'h0D1A: d <= 8'hC0; 15'h0D1B: d <= 8'hC0;
                15'h0D1C: d <= 8'hC0; 15'h0D1D: d <= 8'hC0; 15'h0D1E: d <= 8'hC0; 15'h0D1F: d <= 8'hC0;
                15'h0D20: d <= 8'hC0; 15'h0D21: d <= 8'hC0; 15'h0D22: d <= 8'hC0; 15'h0D23: d <= 8'hC0;
                15'h0D24: d <= 8'hC0; 15'h0D25: d <= 8'hC0; 15'h0D26: d <= 8'hC0; 15'h0D27: d <= 8'hC0;
                15'h0D28: d <= 8'hC0; 15'h0D29: d <= 8'hC0; 15'h0D2A: d <= 8'hC0; 15'h0D2B: d <= 8'hC0;
                15'h0D2C: d <= 8'hC0; 15'h0D2D: d <= 8'hC0; 15'h0D2E: d <= 8'hC0; 15'h0D2F: d <= 8'hC0;
                15'h0D30: d <= 8'hC0; 15'h0D31: d <= 8'hC0; 15'h0D32: d <= 8'hC0; 15'h0D33: d <= 8'hC0;
                15'h0D34: d <= 8'hC0; 15'h0D35: d <= 8'hC0; 15'h0D36: d <= 8'hC0; 15'h0D37: d <= 8'hC0;
                15'h0D38: d <= 8'hC0; 15'h0D39: d <= 8'hC0; 15'h0D3A: d <= 8'hC0; 15'h0D3B: d <= 8'hC0;
                15'h0D3C: d <= 8'hC0; 15'h0D3D: d <= 8'hC0; 15'h0D3E: d <= 8'hC0; 15'h0D3F: d <= 8'hC0;
                15'h0D40: d <= 8'hC0; 15'h0D41: d <= 8'hC0; 15'h0D42: d <= 8'hC0; 15'h0D43: d <= 8'hC0;
                15'h0D44: d <= 8'hC0; 15'h0D45: d <= 8'hC0; 15'h0D46: d <= 8'hC0; 15'h0D47: d <= 8'hC0;
                15'h0D48: d <= 8'hC0; 15'h0D49: d <= 8'hC0; 15'h0D4A: d <= 8'hC0; 15'h0D4B: d <= 8'hC0;
                15'h0D4C: d <= 8'hC0; 15'h0D4D: d <= 8'hC0; 15'h0D4E: d <= 8'hC0; 15'h0D4F: d <= 8'hC0;
                15'h0D50: d <= 8'hC0; 15'h0D51: d <= 8'hC0; 15'h0D52: d <= 8'hC0; 15'h0D53: d <= 8'hC0;
                15'h0D54: d <= 8'hC0; 15'h0D55: d <= 8'hC0; 15'h0D56: d <= 8'hC0; 15'h0D57: d <= 8'hC0;
                15'h0D58: d <= 8'hC0; 15'h0D59: d <= 8'hC0; 15'h0D5A: d <= 8'hC0; 15'h0D5B: d <= 8'hC0;
                15'h0D5C: d <= 8'hC0; 15'h0D5D: d <= 8'hC0; 15'h0D5E: d <= 8'hC0; 15'h0D5F: d <= 8'hC0;
                15'h0D60: d <= 8'hC0; 15'h0D61: d <= 8'hC0; 15'h0D62: d <= 8'hC0; 15'h0D63: d <= 8'hC0;
                15'h0D64: d <= 8'hC0; 15'h0D65: d <= 8'hC0; 15'h0D66: d <= 8'hC0; 15'h0D67: d <= 8'hC0;
                15'h0D68: d <= 8'hC0; 15'h0D69: d <= 8'hC0; 15'h0D6A: d <= 8'hC0; 15'h0D6B: d <= 8'hC0;
                15'h0D6C: d <= 8'hC0; 15'h0D6D: d <= 8'hC0; 15'h0D6E: d <= 8'hC0; 15'h0D6F: d <= 8'hC0;
                15'h0D70: d <= 8'hC0; 15'h0D71: d <= 8'hC0; 15'h0D72: d <= 8'hC0; 15'h0D73: d <= 8'hC0;
                15'h0D74: d <= 8'hC0; 15'h0D75: d <= 8'hC0; 15'h0D76: d <= 8'hC0; 15'h0D77: d <= 8'hC0;
                15'h0D78: d <= 8'hC0; 15'h0D79: d <= 8'hC0; 15'h0D7A: d <= 8'hC0; 15'h0D7B: d <= 8'hC0;
                15'h0D7C: d <= 8'hC0; 15'h0D7D: d <= 8'hC0; 15'h0D7E: d <= 8'hC0; 15'h0D7F: d <= 8'hC0;
                15'h0D80: d <= 8'hC0; 15'h0D81: d <= 8'hC0; 15'h0D82: d <= 8'hC0; 15'h0D83: d <= 8'hC0;
                15'h0D84: d <= 8'hC0; 15'h0D85: d <= 8'hC0; 15'h0D86: d <= 8'hC0; 15'h0D87: d <= 8'hC0;
                15'h0D88: d <= 8'hC0; 15'h0D89: d <= 8'hC0; 15'h0D8A: d <= 8'hC0; 15'h0D8B: d <= 8'hC0;
                15'h0D8C: d <= 8'hC0; 15'h0D8D: d <= 8'hC0; 15'h0D8E: d <= 8'hC0; 15'h0D8F: d <= 8'hC0;
                15'h0D90: d <= 8'hC0; 15'h0D91: d <= 8'hC0; 15'h0D92: d <= 8'hC0; 15'h0D93: d <= 8'hC0;
                15'h0D94: d <= 8'hC0; 15'h0D95: d <= 8'hC0; 15'h0D96: d <= 8'hC0; 15'h0D97: d <= 8'hC0;
                15'h0D98: d <= 8'hC0; 15'h0D99: d <= 8'hC0; 15'h0D9A: d <= 8'hC0; 15'h0D9B: d <= 8'hC0;
                15'h0D9C: d <= 8'hC0; 15'h0D9D: d <= 8'hC0; 15'h0D9E: d <= 8'hC0; 15'h0D9F: d <= 8'hC0;
                15'h0DA0: d <= 8'hC0; 15'h0DA1: d <= 8'hC0; 15'h0DA2: d <= 8'hC0; 15'h0DA3: d <= 8'hC0;
                15'h0DA4: d <= 8'hC0; 15'h0DA5: d <= 8'hC0; 15'h0DA6: d <= 8'hC0; 15'h0DA7: d <= 8'hC0;
                15'h0DA8: d <= 8'hC0; 15'h0DA9: d <= 8'hC0; 15'h0DAA: d <= 8'hC0; 15'h0DAB: d <= 8'hC0;
                15'h0DAC: d <= 8'hC0; 15'h0DAD: d <= 8'hC0; 15'h0DAE: d <= 8'hC0; 15'h0DAF: d <= 8'hC0;
                15'h0DB0: d <= 8'hC0; 15'h0DB1: d <= 8'hC0; 15'h0DB2: d <= 8'hC0; 15'h0DB3: d <= 8'hC0;
                15'h0DB4: d <= 8'hC0; 15'h0DB5: d <= 8'hC0; 15'h0DB6: d <= 8'hC0; 15'h0DB7: d <= 8'hC0;
                15'h0DB8: d <= 8'hC0; 15'h0DB9: d <= 8'hC0; 15'h0DBA: d <= 8'hC0; 15'h0DBB: d <= 8'hC0;
                15'h0DBC: d <= 8'hC0; 15'h0DBD: d <= 8'hC0; 15'h0DBE: d <= 8'hC0; 15'h0DBF: d <= 8'hC0;
                15'h0DC0: d <= 8'hC0; 15'h0DC1: d <= 8'hC0; 15'h0DC2: d <= 8'hC0; 15'h0DC3: d <= 8'hC0;
                15'h0DC4: d <= 8'hC0; 15'h0DC5: d <= 8'hC0; 15'h0DC6: d <= 8'hC0; 15'h0DC7: d <= 8'hC0;
                15'h0DC8: d <= 8'hC0; 15'h0DC9: d <= 8'hC0; 15'h0DCA: d <= 8'hC0; 15'h0DCB: d <= 8'hC0;
                15'h0DCC: d <= 8'hC0; 15'h0DCD: d <= 8'hC0; 15'h0DCE: d <= 8'hC0; 15'h0DCF: d <= 8'hC0;
                15'h0DD0: d <= 8'hC0; 15'h0DD1: d <= 8'hC0; 15'h0DD2: d <= 8'hC0; 15'h0DD3: d <= 8'hC0;
                15'h0DD4: d <= 8'hC0; 15'h0DD5: d <= 8'hC0; 15'h0DD6: d <= 8'hC0; 15'h0DD7: d <= 8'hC0;
                15'h0DD8: d <= 8'hC0; 15'h0DD9: d <= 8'hC0; 15'h0DDA: d <= 8'hC0; 15'h0DDB: d <= 8'hC0;
                15'h0DDC: d <= 8'hC0; 15'h0DDD: d <= 8'hC0; 15'h0DDE: d <= 8'hC0; 15'h0DDF: d <= 8'hC0;
                15'h0DE0: d <= 8'hC0; 15'h0DE1: d <= 8'hC0; 15'h0DE2: d <= 8'hC0; 15'h0DE3: d <= 8'hC0;
                15'h0DE4: d <= 8'hC0; 15'h0DE5: d <= 8'hC0; 15'h0DE6: d <= 8'hC0; 15'h0DE7: d <= 8'hC0;
                15'h0DE8: d <= 8'hC0; 15'h0DE9: d <= 8'hC0; 15'h0DEA: d <= 8'hC0; 15'h0DEB: d <= 8'hC0;
                15'h0DEC: d <= 8'hC0; 15'h0DED: d <= 8'hC0; 15'h0DEE: d <= 8'hC0; 15'h0DEF: d <= 8'hC0;
                15'h0DF0: d <= 8'hC0; 15'h0DF1: d <= 8'hC0; 15'h0DF2: d <= 8'hC0; 15'h0DF3: d <= 8'hC0;
                15'h0DF4: d <= 8'hC0; 15'h0DF5: d <= 8'hC0; 15'h0DF6: d <= 8'hC0; 15'h0DF7: d <= 8'hC0;
                15'h0DF8: d <= 8'hC0; 15'h0DF9: d <= 8'hC0; 15'h0DFA: d <= 8'hC0; 15'h0DFB: d <= 8'hC0;
                15'h0DFC: d <= 8'hC0; 15'h0DFD: d <= 8'hC0; 15'h0DFE: d <= 8'hC0; 15'h0DFF: d <= 8'hC0;
                15'h0E00: d <= 8'hC0; 15'h0E01: d <= 8'hC0; 15'h0E02: d <= 8'hC0; 15'h0E03: d <= 8'hC0;
                15'h0E04: d <= 8'hC0; 15'h0E05: d <= 8'hC0; 15'h0E06: d <= 8'hC0; 15'h0E07: d <= 8'hC0;
                15'h0E08: d <= 8'hC0; 15'h0E09: d <= 8'hC0; 15'h0E0A: d <= 8'hC0; 15'h0E0B: d <= 8'hC0;
                15'h0E0C: d <= 8'hC0; 15'h0E0D: d <= 8'hC0; 15'h0E0E: d <= 8'hC0; 15'h0E0F: d <= 8'hC0;
                15'h0E10: d <= 8'hC0; 15'h0E11: d <= 8'hC0; 15'h0E12: d <= 8'hC0; 15'h0E13: d <= 8'hC0;
                15'h0E14: d <= 8'hC0; 15'h0E15: d <= 8'hC0; 15'h0E16: d <= 8'hC0; 15'h0E17: d <= 8'hC0;
                15'h0E18: d <= 8'hC0; 15'h0E19: d <= 8'hC0; 15'h0E1A: d <= 8'hC0; 15'h0E1B: d <= 8'hC0;
                15'h0E1C: d <= 8'hC0; 15'h0E1D: d <= 8'hC0; 15'h0E1E: d <= 8'hC0; 15'h0E1F: d <= 8'hC0;
                15'h0E20: d <= 8'hC0; 15'h0E21: d <= 8'hC0; 15'h0E22: d <= 8'hC0; 15'h0E23: d <= 8'hC0;
                15'h0E24: d <= 8'hC0; 15'h0E25: d <= 8'hC0; 15'h0E26: d <= 8'hC0; 15'h0E27: d <= 8'hC0;
                15'h0E28: d <= 8'hC0; 15'h0E29: d <= 8'hC0; 15'h0E2A: d <= 8'hC0; 15'h0E2B: d <= 8'hC0;
                15'h0E2C: d <= 8'hC0; 15'h0E2D: d <= 8'hC0; 15'h0E2E: d <= 8'hC0; 15'h0E2F: d <= 8'hC0;
                15'h0E30: d <= 8'hC0; 15'h0E31: d <= 8'hC0; 15'h0E32: d <= 8'hC0; 15'h0E33: d <= 8'hC0;
                15'h0E34: d <= 8'hC0; 15'h0E35: d <= 8'hC0; 15'h0E36: d <= 8'hC0; 15'h0E37: d <= 8'hC0;
                15'h0E38: d <= 8'hC0; 15'h0E39: d <= 8'hC0; 15'h0E3A: d <= 8'hC0; 15'h0E3B: d <= 8'hC0;
                15'h0E3C: d <= 8'hC0; 15'h0E3D: d <= 8'hC0; 15'h0E3E: d <= 8'hC0; 15'h0E3F: d <= 8'hC0;
                15'h0E40: d <= 8'hC0; 15'h0E41: d <= 8'hC0; 15'h0E42: d <= 8'hC0; 15'h0E43: d <= 8'hC0;
                15'h0E44: d <= 8'hC0; 15'h0E45: d <= 8'hC0; 15'h0E46: d <= 8'hC0; 15'h0E47: d <= 8'hC0;
                15'h0E48: d <= 8'hC0; 15'h0E49: d <= 8'hC0; 15'h0E4A: d <= 8'hC0; 15'h0E4B: d <= 8'hC0;
                15'h0E4C: d <= 8'hC0; 15'h0E4D: d <= 8'hC0; 15'h0E4E: d <= 8'hC0; 15'h0E4F: d <= 8'hC0;
                15'h0E50: d <= 8'hC0; 15'h0E51: d <= 8'hC0; 15'h0E52: d <= 8'hC0; 15'h0E53: d <= 8'hC0;
                15'h0E54: d <= 8'hC0; 15'h0E55: d <= 8'hC0; 15'h0E56: d <= 8'hC0; 15'h0E57: d <= 8'hC0;
                15'h0E58: d <= 8'hC0; 15'h0E59: d <= 8'hC0; 15'h0E5A: d <= 8'hC0; 15'h0E5B: d <= 8'hC0;
                15'h0E5C: d <= 8'hC0; 15'h0E5D: d <= 8'hC0; 15'h0E5E: d <= 8'hC0; 15'h0E5F: d <= 8'hC0;
                15'h0E60: d <= 8'hC0; 15'h0E61: d <= 8'hC0; 15'h0E62: d <= 8'hC0; 15'h0E63: d <= 8'hC0;
                15'h0E64: d <= 8'hC0; 15'h0E65: d <= 8'hC0; 15'h0E66: d <= 8'hC0; 15'h0E67: d <= 8'hC0;
                15'h0E68: d <= 8'hC0; 15'h0E69: d <= 8'hC0; 15'h0E6A: d <= 8'hC0; 15'h0E6B: d <= 8'hC0;
                15'h0E6C: d <= 8'hC0; 15'h0E6D: d <= 8'hC0; 15'h0E6E: d <= 8'hC0; 15'h0E6F: d <= 8'hC0;
                15'h0E70: d <= 8'hC0; 15'h0E71: d <= 8'hC0; 15'h0E72: d <= 8'hC0; 15'h0E73: d <= 8'hC0;
                15'h0E74: d <= 8'hC0; 15'h0E75: d <= 8'hC0; 15'h0E76: d <= 8'hC0; 15'h0E77: d <= 8'hC0;
                15'h0E78: d <= 8'hC0; 15'h0E79: d <= 8'hC0; 15'h0E7A: d <= 8'hC0; 15'h0E7B: d <= 8'hC0;
                15'h0E7C: d <= 8'hC0; 15'h0E7D: d <= 8'hC0; 15'h0E7E: d <= 8'hC0; 15'h0E7F: d <= 8'hC0;
                15'h0E80: d <= 8'hC0; 15'h0E81: d <= 8'hC0; 15'h0E82: d <= 8'hC0; 15'h0E83: d <= 8'hC0;
                15'h0E84: d <= 8'hC0; 15'h0E85: d <= 8'hC0; 15'h0E86: d <= 8'hC0; 15'h0E87: d <= 8'hC0;
                15'h0E88: d <= 8'hC0; 15'h0E89: d <= 8'hC0; 15'h0E8A: d <= 8'hC0; 15'h0E8B: d <= 8'hC0;
                15'h0E8C: d <= 8'hC0; 15'h0E8D: d <= 8'hC0; 15'h0E8E: d <= 8'hC0; 15'h0E8F: d <= 8'hC0;
                15'h0E90: d <= 8'hC0; 15'h0E91: d <= 8'hC0; 15'h0E92: d <= 8'hC0; 15'h0E93: d <= 8'hC0;
                15'h0E94: d <= 8'hC0; 15'h0E95: d <= 8'hC0; 15'h0E96: d <= 8'hC0; 15'h0E97: d <= 8'hC0;
                15'h0E98: d <= 8'hC0; 15'h0E99: d <= 8'hC0; 15'h0E9A: d <= 8'hC0; 15'h0E9B: d <= 8'hC0;
                15'h0E9C: d <= 8'hC0; 15'h0E9D: d <= 8'hC0; 15'h0E9E: d <= 8'hC0; 15'h0E9F: d <= 8'hC0;
                15'h0EA0: d <= 8'hC0; 15'h0EA1: d <= 8'hC0; 15'h0EA2: d <= 8'hC0; 15'h0EA3: d <= 8'hC0;
                15'h0EA4: d <= 8'hC0; 15'h0EA5: d <= 8'hC0; 15'h0EA6: d <= 8'hC0; 15'h0EA7: d <= 8'hC0;
                15'h0EA8: d <= 8'hC0; 15'h0EA9: d <= 8'hC0; 15'h0EAA: d <= 8'hC0; 15'h0EAB: d <= 8'hC0;
                15'h0EAC: d <= 8'hC0; 15'h0EAD: d <= 8'hC0; 15'h0EAE: d <= 8'hC0; 15'h0EAF: d <= 8'hC0;
                15'h0EB0: d <= 8'hC0; 15'h0EB1: d <= 8'hC0; 15'h0EB2: d <= 8'hC0; 15'h0EB3: d <= 8'hC0;
                15'h0EB4: d <= 8'hC0; 15'h0EB5: d <= 8'hC0; 15'h0EB6: d <= 8'hC0; 15'h0EB7: d <= 8'hC0;
                15'h0EB8: d <= 8'hC0; 15'h0EB9: d <= 8'hC0; 15'h0EBA: d <= 8'hC0; 15'h0EBB: d <= 8'hC0;
                15'h0EBC: d <= 8'hC0; 15'h0EBD: d <= 8'hC0; 15'h0EBE: d <= 8'hC0; 15'h0EBF: d <= 8'hC0;
                15'h0EC0: d <= 8'hC0; 15'h0EC1: d <= 8'hC0; 15'h0EC2: d <= 8'hC0; 15'h0EC3: d <= 8'hC0;
                15'h0EC4: d <= 8'hC0; 15'h0EC5: d <= 8'hC0; 15'h0EC6: d <= 8'hC0; 15'h0EC7: d <= 8'hC0;
                15'h0EC8: d <= 8'hC0; 15'h0EC9: d <= 8'hC0; 15'h0ECA: d <= 8'hC0; 15'h0ECB: d <= 8'hC0;
                15'h0ECC: d <= 8'hC0; 15'h0ECD: d <= 8'hC0; 15'h0ECE: d <= 8'hC0; 15'h0ECF: d <= 8'hC0;
                15'h0ED0: d <= 8'hC0; 15'h0ED1: d <= 8'hC0; 15'h0ED2: d <= 8'hC0; 15'h0ED3: d <= 8'hC0;
                15'h0ED4: d <= 8'hC0; 15'h0ED5: d <= 8'hC0; 15'h0ED6: d <= 8'hC0; 15'h0ED7: d <= 8'hC0;
                15'h0ED8: d <= 8'hC0; 15'h0ED9: d <= 8'hC0; 15'h0EDA: d <= 8'hC0; 15'h0EDB: d <= 8'hC0;
                15'h0EDC: d <= 8'hC0; 15'h0EDD: d <= 8'hC0; 15'h0EDE: d <= 8'hC0; 15'h0EDF: d <= 8'hC0;
                15'h0EE0: d <= 8'hC0; 15'h0EE1: d <= 8'hC0; 15'h0EE2: d <= 8'hC0; 15'h0EE3: d <= 8'hC0;
                15'h0EE4: d <= 8'hC0; 15'h0EE5: d <= 8'hC0; 15'h0EE6: d <= 8'hC0; 15'h0EE7: d <= 8'hC0;
                15'h0EE8: d <= 8'hC0; 15'h0EE9: d <= 8'hC0; 15'h0EEA: d <= 8'hC0; 15'h0EEB: d <= 8'hC0;
                15'h0EEC: d <= 8'hC0; 15'h0EED: d <= 8'hC0; 15'h0EEE: d <= 8'hC0; 15'h0EEF: d <= 8'hC0;
                15'h0EF0: d <= 8'hC0; 15'h0EF1: d <= 8'hC0; 15'h0EF2: d <= 8'hC0; 15'h0EF3: d <= 8'hC0;
                15'h0EF4: d <= 8'hC0; 15'h0EF5: d <= 8'hC0; 15'h0EF6: d <= 8'hC0; 15'h0EF7: d <= 8'hC0;
                15'h0EF8: d <= 8'hC0; 15'h0EF9: d <= 8'hC0; 15'h0EFA: d <= 8'hC0; 15'h0EFB: d <= 8'hC0;
                15'h0EFC: d <= 8'hC0; 15'h0EFD: d <= 8'hC0; 15'h0EFE: d <= 8'hC0; 15'h0EFF: d <= 8'hC0;
                15'h0F00: d <= 8'hC0; 15'h0F01: d <= 8'hC0; 15'h0F02: d <= 8'hC0; 15'h0F03: d <= 8'hC0;
                15'h0F04: d <= 8'hC0; 15'h0F05: d <= 8'hC0; 15'h0F06: d <= 8'hC0; 15'h0F07: d <= 8'hC0;
                15'h0F08: d <= 8'hC0; 15'h0F09: d <= 8'hC0; 15'h0F0A: d <= 8'hC0; 15'h0F0B: d <= 8'hC0;
                15'h0F0C: d <= 8'hC0; 15'h0F0D: d <= 8'hC0; 15'h0F0E: d <= 8'hC0; 15'h0F0F: d <= 8'hC0;
                15'h0F10: d <= 8'hC0; 15'h0F11: d <= 8'hC0; 15'h0F12: d <= 8'hC0; 15'h0F13: d <= 8'hC0;
                15'h0F14: d <= 8'hC0; 15'h0F15: d <= 8'hC0; 15'h0F16: d <= 8'hC0; 15'h0F17: d <= 8'hC0;
                15'h0F18: d <= 8'hC0; 15'h0F19: d <= 8'hC0; 15'h0F1A: d <= 8'hC0; 15'h0F1B: d <= 8'hC0;
                15'h0F1C: d <= 8'hC0; 15'h0F1D: d <= 8'hC0; 15'h0F1E: d <= 8'hC0; 15'h0F1F: d <= 8'hC0;
                15'h0F20: d <= 8'hC0; 15'h0F21: d <= 8'hC0; 15'h0F22: d <= 8'hC0; 15'h0F23: d <= 8'hC0;
                15'h0F24: d <= 8'hC0; 15'h0F25: d <= 8'hC0; 15'h0F26: d <= 8'hC0; 15'h0F27: d <= 8'hC0;
                15'h0F28: d <= 8'hC0; 15'h0F29: d <= 8'hC0; 15'h0F2A: d <= 8'hC0; 15'h0F2B: d <= 8'hC0;
                15'h0F2C: d <= 8'hC0; 15'h0F2D: d <= 8'hC0; 15'h0F2E: d <= 8'hC0; 15'h0F2F: d <= 8'hC0;
                15'h0F30: d <= 8'hC0; 15'h0F31: d <= 8'hC0; 15'h0F32: d <= 8'hC0; 15'h0F33: d <= 8'hC0;
                15'h0F34: d <= 8'hC0; 15'h0F35: d <= 8'hC0; 15'h0F36: d <= 8'hC0; 15'h0F37: d <= 8'hC0;
                15'h0F38: d <= 8'hC0; 15'h0F39: d <= 8'hC0; 15'h0F3A: d <= 8'hC0; 15'h0F3B: d <= 8'hC0;
                15'h0F3C: d <= 8'hC0; 15'h0F3D: d <= 8'hC0; 15'h0F3E: d <= 8'hC0; 15'h0F3F: d <= 8'hC0;
                15'h0F40: d <= 8'hC0; 15'h0F41: d <= 8'hC0; 15'h0F42: d <= 8'hC0; 15'h0F43: d <= 8'hC0;
                15'h0F44: d <= 8'hC0; 15'h0F45: d <= 8'hC0; 15'h0F46: d <= 8'hC0; 15'h0F47: d <= 8'hC0;
                15'h0F48: d <= 8'hC0; 15'h0F49: d <= 8'hC0; 15'h0F4A: d <= 8'hC0; 15'h0F4B: d <= 8'hC0;
                15'h0F4C: d <= 8'hC0; 15'h0F4D: d <= 8'hC0; 15'h0F4E: d <= 8'hC0; 15'h0F4F: d <= 8'hC0;
                15'h0F50: d <= 8'hC0; 15'h0F51: d <= 8'hC0; 15'h0F52: d <= 8'hC0; 15'h0F53: d <= 8'hC0;
                15'h0F54: d <= 8'hC0; 15'h0F55: d <= 8'hC0; 15'h0F56: d <= 8'hC0; 15'h0F57: d <= 8'hC0;
                15'h0F58: d <= 8'hC0; 15'h0F59: d <= 8'hC0; 15'h0F5A: d <= 8'hC0; 15'h0F5B: d <= 8'hC0;
                15'h0F5C: d <= 8'hC0; 15'h0F5D: d <= 8'hC0; 15'h0F5E: d <= 8'hC0; 15'h0F5F: d <= 8'hC0;
                15'h0F60: d <= 8'hC0; 15'h0F61: d <= 8'hC0; 15'h0F62: d <= 8'hC0; 15'h0F63: d <= 8'hC0;
                15'h0F64: d <= 8'hC0; 15'h0F65: d <= 8'hC0; 15'h0F66: d <= 8'hC0; 15'h0F67: d <= 8'hC0;
                15'h0F68: d <= 8'hC0; 15'h0F69: d <= 8'hC0; 15'h0F6A: d <= 8'hC0; 15'h0F6B: d <= 8'hC0;
                15'h0F6C: d <= 8'hC0; 15'h0F6D: d <= 8'hC0; 15'h0F6E: d <= 8'hC0; 15'h0F6F: d <= 8'hC0;
                15'h0F70: d <= 8'hC0; 15'h0F71: d <= 8'hC0; 15'h0F72: d <= 8'hC0; 15'h0F73: d <= 8'hC0;
                15'h0F74: d <= 8'hC0; 15'h0F75: d <= 8'hC0; 15'h0F76: d <= 8'hC0; 15'h0F77: d <= 8'hC0;
                15'h0F78: d <= 8'hC0; 15'h0F79: d <= 8'hC0; 15'h0F7A: d <= 8'hC0; 15'h0F7B: d <= 8'hC0;
                15'h0F7C: d <= 8'hC0; 15'h0F7D: d <= 8'hC0; 15'h0F7E: d <= 8'hC0; 15'h0F7F: d <= 8'hC0;
                15'h0F80: d <= 8'hC0; 15'h0F81: d <= 8'hC0; 15'h0F82: d <= 8'hC0; 15'h0F83: d <= 8'hC0;
                15'h0F84: d <= 8'hC0; 15'h0F85: d <= 8'hC0; 15'h0F86: d <= 8'hC0; 15'h0F87: d <= 8'hC0;
                15'h0F88: d <= 8'hC0; 15'h0F89: d <= 8'hC0; 15'h0F8A: d <= 8'hC0; 15'h0F8B: d <= 8'hC0;
                15'h0F8C: d <= 8'hC0; 15'h0F8D: d <= 8'hC0; 15'h0F8E: d <= 8'hC0; 15'h0F8F: d <= 8'hC0;
                15'h0F90: d <= 8'hC0; 15'h0F91: d <= 8'hC0; 15'h0F92: d <= 8'hC0; 15'h0F93: d <= 8'hC0;
                15'h0F94: d <= 8'hC0; 15'h0F95: d <= 8'hC0; 15'h0F96: d <= 8'hC0; 15'h0F97: d <= 8'hC0;
                15'h0F98: d <= 8'hC0; 15'h0F99: d <= 8'hC0; 15'h0F9A: d <= 8'hC0; 15'h0F9B: d <= 8'hC0;
                15'h0F9C: d <= 8'hC0; 15'h0F9D: d <= 8'hC0; 15'h0F9E: d <= 8'hC0; 15'h0F9F: d <= 8'hC0;
                15'h0FA0: d <= 8'hC0; 15'h0FA1: d <= 8'hC0; 15'h0FA2: d <= 8'hC0; 15'h0FA3: d <= 8'hC0;
                15'h0FA4: d <= 8'hC0; 15'h0FA5: d <= 8'hC0; 15'h0FA6: d <= 8'hC0; 15'h0FA7: d <= 8'hC0;
                15'h0FA8: d <= 8'hC0; 15'h0FA9: d <= 8'hC0; 15'h0FAA: d <= 8'hC0; 15'h0FAB: d <= 8'hC0;
                15'h0FAC: d <= 8'hC0; 15'h0FAD: d <= 8'hC0; 15'h0FAE: d <= 8'hC0; 15'h0FAF: d <= 8'hC0;
                15'h0FB0: d <= 8'hC0; 15'h0FB1: d <= 8'hC0; 15'h0FB2: d <= 8'hC0; 15'h0FB3: d <= 8'hC0;
                15'h0FB4: d <= 8'hC0; 15'h0FB5: d <= 8'hC0; 15'h0FB6: d <= 8'hC0; 15'h0FB7: d <= 8'hC0;
                15'h0FB8: d <= 8'hC0; 15'h0FB9: d <= 8'hC0; 15'h0FBA: d <= 8'hC0; 15'h0FBB: d <= 8'hC0;
                15'h0FBC: d <= 8'hC0; 15'h0FBD: d <= 8'hC0; 15'h0FBE: d <= 8'hC0; 15'h0FBF: d <= 8'hC0;
                15'h0FC0: d <= 8'hC0; 15'h0FC1: d <= 8'hC0; 15'h0FC2: d <= 8'hC0; 15'h0FC3: d <= 8'hC0;
                15'h0FC4: d <= 8'hC0; 15'h0FC5: d <= 8'hC0; 15'h0FC6: d <= 8'hC0; 15'h0FC7: d <= 8'hC0;
                15'h0FC8: d <= 8'hC0; 15'h0FC9: d <= 8'hC0; 15'h0FCA: d <= 8'hC0; 15'h0FCB: d <= 8'hC0;
                15'h0FCC: d <= 8'hC0; 15'h0FCD: d <= 8'hC0; 15'h0FCE: d <= 8'hC0; 15'h0FCF: d <= 8'hC0;
                15'h0FD0: d <= 8'hC0; 15'h0FD1: d <= 8'hC0; 15'h0FD2: d <= 8'hC0; 15'h0FD3: d <= 8'hC0;
                15'h0FD4: d <= 8'hC0; 15'h0FD5: d <= 8'hC0; 15'h0FD6: d <= 8'hC0; 15'h0FD7: d <= 8'hC0;
                15'h0FD8: d <= 8'hC0; 15'h0FD9: d <= 8'hC0; 15'h0FDA: d <= 8'hC0; 15'h0FDB: d <= 8'hC0;
                15'h0FDC: d <= 8'hC0; 15'h0FDD: d <= 8'hC0; 15'h0FDE: d <= 8'hC0; 15'h0FDF: d <= 8'hC0;
                15'h0FE0: d <= 8'hC0; 15'h0FE1: d <= 8'hC0; 15'h0FE2: d <= 8'hC0; 15'h0FE3: d <= 8'hC0;
                15'h0FE4: d <= 8'hC0; 15'h0FE5: d <= 8'hC0; 15'h0FE6: d <= 8'hC0; 15'h0FE7: d <= 8'hC0;
                15'h0FE8: d <= 8'hC0; 15'h0FE9: d <= 8'hC0; 15'h0FEA: d <= 8'hC0; 15'h0FEB: d <= 8'hC0;
                15'h0FEC: d <= 8'hC0; 15'h0FED: d <= 8'hC0; 15'h0FEE: d <= 8'hC0; 15'h0FEF: d <= 8'hC0;
                15'h0FF0: d <= 8'hC0; 15'h0FF1: d <= 8'hC0; 15'h0FF2: d <= 8'hC0; 15'h0FF3: d <= 8'hC0;
                15'h0FF4: d <= 8'hC0; 15'h0FF5: d <= 8'hC0; 15'h0FF6: d <= 8'hC0; 15'h0FF7: d <= 8'hC0;
                15'h0FF8: d <= 8'hC0; 15'h0FF9: d <= 8'hC0; 15'h0FFA: d <= 8'hC0; 15'h0FFB: d <= 8'hC0;
                15'h0FFC: d <= 8'hC0; 15'h0FFD: d <= 8'hC0; 15'h0FFE: d <= 8'hC0; 15'h0FFF: d <= 8'hC0;
                15'h1000: d <= 8'hC0; 15'h1001: d <= 8'hC0; 15'h1002: d <= 8'hC0; 15'h1003: d <= 8'hC0;
                15'h1004: d <= 8'hC0; 15'h1005: d <= 8'hC0; 15'h1006: d <= 8'hC0; 15'h1007: d <= 8'hC0;
                15'h1008: d <= 8'hC0; 15'h1009: d <= 8'hC0; 15'h100A: d <= 8'hC0; 15'h100B: d <= 8'hC0;
                15'h100C: d <= 8'hC0; 15'h100D: d <= 8'hC0; 15'h100E: d <= 8'hC0; 15'h100F: d <= 8'hC0;
                15'h1010: d <= 8'hC0; 15'h1011: d <= 8'hC0; 15'h1012: d <= 8'hC0; 15'h1013: d <= 8'hC0;
                15'h1014: d <= 8'hC0; 15'h1015: d <= 8'hC0; 15'h1016: d <= 8'hC0; 15'h1017: d <= 8'hC0;
                15'h1018: d <= 8'hC0; 15'h1019: d <= 8'hC0; 15'h101A: d <= 8'hC0; 15'h101B: d <= 8'hC0;
                15'h101C: d <= 8'hC0; 15'h101D: d <= 8'hC0; 15'h101E: d <= 8'hC0; 15'h101F: d <= 8'hC0;
                15'h1020: d <= 8'hC0; 15'h1021: d <= 8'hC0; 15'h1022: d <= 8'hC0; 15'h1023: d <= 8'hC0;
                15'h1024: d <= 8'hC0; 15'h1025: d <= 8'hC0; 15'h1026: d <= 8'hC0; 15'h1027: d <= 8'hC0;
                15'h1028: d <= 8'hC0; 15'h1029: d <= 8'hC0; 15'h102A: d <= 8'hC0; 15'h102B: d <= 8'hC0;
                15'h102C: d <= 8'hC0; 15'h102D: d <= 8'hC0; 15'h102E: d <= 8'hC0; 15'h102F: d <= 8'hC0;
                15'h1030: d <= 8'hC0; 15'h1031: d <= 8'hC0; 15'h1032: d <= 8'hC0; 15'h1033: d <= 8'hC0;
                15'h1034: d <= 8'hC0; 15'h1035: d <= 8'hC0; 15'h1036: d <= 8'hC0; 15'h1037: d <= 8'hC0;
                15'h1038: d <= 8'hC0; 15'h1039: d <= 8'hC0; 15'h103A: d <= 8'hC0; 15'h103B: d <= 8'hC0;
                15'h103C: d <= 8'hC0; 15'h103D: d <= 8'hC0; 15'h103E: d <= 8'hC0; 15'h103F: d <= 8'hC0;
                15'h1040: d <= 8'hC0; 15'h1041: d <= 8'hC0; 15'h1042: d <= 8'hC0; 15'h1043: d <= 8'hC0;
                15'h1044: d <= 8'hC0; 15'h1045: d <= 8'hC0; 15'h1046: d <= 8'hC0; 15'h1047: d <= 8'hC0;
                15'h1048: d <= 8'hC0; 15'h1049: d <= 8'hC0; 15'h104A: d <= 8'hC0; 15'h104B: d <= 8'hC0;
                15'h104C: d <= 8'hC0; 15'h104D: d <= 8'hC0; 15'h104E: d <= 8'hC0; 15'h104F: d <= 8'hC0;
                15'h1050: d <= 8'hC0; 15'h1051: d <= 8'hC0; 15'h1052: d <= 8'hC0; 15'h1053: d <= 8'hC0;
                15'h1054: d <= 8'hC0; 15'h1055: d <= 8'hC0; 15'h1056: d <= 8'hC0; 15'h1057: d <= 8'hC0;
                15'h1058: d <= 8'hC0; 15'h1059: d <= 8'hC0; 15'h105A: d <= 8'hC0; 15'h105B: d <= 8'hC0;
                15'h105C: d <= 8'hC0; 15'h105D: d <= 8'hC0; 15'h105E: d <= 8'hC0; 15'h105F: d <= 8'hC0;
                15'h1060: d <= 8'hC0; 15'h1061: d <= 8'hC0; 15'h1062: d <= 8'hC0; 15'h1063: d <= 8'hC0;
                15'h1064: d <= 8'hC0; 15'h1065: d <= 8'hC0; 15'h1066: d <= 8'hC0; 15'h1067: d <= 8'hC0;
                15'h1068: d <= 8'hC0; 15'h1069: d <= 8'hC0; 15'h106A: d <= 8'hC0; 15'h106B: d <= 8'hC0;
                15'h106C: d <= 8'hC0; 15'h106D: d <= 8'hC0; 15'h106E: d <= 8'hC0; 15'h106F: d <= 8'hC0;
                15'h1070: d <= 8'hC0; 15'h1071: d <= 8'hC0; 15'h1072: d <= 8'hC0; 15'h1073: d <= 8'hC0;
                15'h1074: d <= 8'hC0; 15'h1075: d <= 8'hC0; 15'h1076: d <= 8'hC0; 15'h1077: d <= 8'hC0;
                15'h1078: d <= 8'hC0; 15'h1079: d <= 8'hC0; 15'h107A: d <= 8'hC0; 15'h107B: d <= 8'hC0;
                15'h107C: d <= 8'hC0; 15'h107D: d <= 8'hC0; 15'h107E: d <= 8'hC0; 15'h107F: d <= 8'hC0;
                15'h1080: d <= 8'hC0; 15'h1081: d <= 8'hC0; 15'h1082: d <= 8'hC0; 15'h1083: d <= 8'hC0;
                15'h1084: d <= 8'hC0; 15'h1085: d <= 8'hC0; 15'h1086: d <= 8'hC0; 15'h1087: d <= 8'hC0;
                15'h1088: d <= 8'hC0; 15'h1089: d <= 8'hC0; 15'h108A: d <= 8'hC0; 15'h108B: d <= 8'hC0;
                15'h108C: d <= 8'hC0; 15'h108D: d <= 8'hC0; 15'h108E: d <= 8'hC0; 15'h108F: d <= 8'hC0;
                15'h1090: d <= 8'hC0; 15'h1091: d <= 8'hC0; 15'h1092: d <= 8'hC0; 15'h1093: d <= 8'hC0;
                15'h1094: d <= 8'hC0; 15'h1095: d <= 8'hC0; 15'h1096: d <= 8'hC0; 15'h1097: d <= 8'hC0;
                15'h1098: d <= 8'hC0; 15'h1099: d <= 8'hC0; 15'h109A: d <= 8'hC0; 15'h109B: d <= 8'hC0;
                15'h109C: d <= 8'hC0; 15'h109D: d <= 8'hC0; 15'h109E: d <= 8'hC0; 15'h109F: d <= 8'hC0;
                15'h10A0: d <= 8'hC0; 15'h10A1: d <= 8'hC0; 15'h10A2: d <= 8'hC0; 15'h10A3: d <= 8'hC0;
                15'h10A4: d <= 8'hC0; 15'h10A5: d <= 8'hC0; 15'h10A6: d <= 8'hC0; 15'h10A7: d <= 8'hC0;
                15'h10A8: d <= 8'hC0; 15'h10A9: d <= 8'hC0; 15'h10AA: d <= 8'hC0; 15'h10AB: d <= 8'hC0;
                15'h10AC: d <= 8'hC0; 15'h10AD: d <= 8'hC0; 15'h10AE: d <= 8'hC0; 15'h10AF: d <= 8'hC0;
                15'h10B0: d <= 8'hC0; 15'h10B1: d <= 8'hC0; 15'h10B2: d <= 8'hC0; 15'h10B3: d <= 8'hC0;
                15'h10B4: d <= 8'hC0; 15'h10B5: d <= 8'hC0; 15'h10B6: d <= 8'hC0; 15'h10B7: d <= 8'hC0;
                15'h10B8: d <= 8'hC0; 15'h10B9: d <= 8'hC0; 15'h10BA: d <= 8'hC0; 15'h10BB: d <= 8'hC0;
                15'h10BC: d <= 8'hC0; 15'h10BD: d <= 8'hC0; 15'h10BE: d <= 8'hC0; 15'h10BF: d <= 8'hC0;
                15'h10C0: d <= 8'hC0; 15'h10C1: d <= 8'hC0; 15'h10C2: d <= 8'hC0; 15'h10C3: d <= 8'hC0;
                15'h10C4: d <= 8'hC0; 15'h10C5: d <= 8'hC0; 15'h10C6: d <= 8'hC0; 15'h10C7: d <= 8'hC0;
                15'h10C8: d <= 8'hC0; 15'h10C9: d <= 8'hC0; 15'h10CA: d <= 8'hC0; 15'h10CB: d <= 8'hC0;
                15'h10CC: d <= 8'hC0; 15'h10CD: d <= 8'hC0; 15'h10CE: d <= 8'hC0; 15'h10CF: d <= 8'hC0;
                15'h10D0: d <= 8'hC0; 15'h10D1: d <= 8'hC0; 15'h10D2: d <= 8'hC0; 15'h10D3: d <= 8'hC0;
                15'h10D4: d <= 8'hC0; 15'h10D5: d <= 8'hC0; 15'h10D6: d <= 8'hC0; 15'h10D7: d <= 8'hC0;
                15'h10D8: d <= 8'hC0; 15'h10D9: d <= 8'hC0; 15'h10DA: d <= 8'hC0; 15'h10DB: d <= 8'hC0;
                15'h10DC: d <= 8'hC0; 15'h10DD: d <= 8'hC0; 15'h10DE: d <= 8'hC0; 15'h10DF: d <= 8'hC0;
                15'h10E0: d <= 8'hC0; 15'h10E1: d <= 8'hC0; 15'h10E2: d <= 8'hC0; 15'h10E3: d <= 8'hC0;
                15'h10E4: d <= 8'hC0; 15'h10E5: d <= 8'hC0; 15'h10E6: d <= 8'hC0; 15'h10E7: d <= 8'hC0;
                15'h10E8: d <= 8'hC0; 15'h10E9: d <= 8'hC0; 15'h10EA: d <= 8'hC0; 15'h10EB: d <= 8'hC0;
                15'h10EC: d <= 8'hC0; 15'h10ED: d <= 8'hC0; 15'h10EE: d <= 8'hC0; 15'h10EF: d <= 8'hC0;
                15'h10F0: d <= 8'hC0; 15'h10F1: d <= 8'hC0; 15'h10F2: d <= 8'hC0; 15'h10F3: d <= 8'hC0;
                15'h10F4: d <= 8'hC0; 15'h10F5: d <= 8'hC0; 15'h10F6: d <= 8'hC0; 15'h10F7: d <= 8'hC0;
                15'h10F8: d <= 8'hC0; 15'h10F9: d <= 8'hC0; 15'h10FA: d <= 8'hC0; 15'h10FB: d <= 8'hC0;
                15'h10FC: d <= 8'hC0; 15'h10FD: d <= 8'hC0; 15'h10FE: d <= 8'hC0; 15'h10FF: d <= 8'hC0;
                15'h1100: d <= 8'hC0; 15'h1101: d <= 8'hC0; 15'h1102: d <= 8'hC0; 15'h1103: d <= 8'hC0;
                15'h1104: d <= 8'hC0; 15'h1105: d <= 8'hC0; 15'h1106: d <= 8'hC0; 15'h1107: d <= 8'hC0;
                15'h1108: d <= 8'hC0; 15'h1109: d <= 8'hC0; 15'h110A: d <= 8'hC0; 15'h110B: d <= 8'hC0;
                15'h110C: d <= 8'hC0; 15'h110D: d <= 8'hC0; 15'h110E: d <= 8'hC0; 15'h110F: d <= 8'hC0;
                15'h1110: d <= 8'hC0; 15'h1111: d <= 8'hC0; 15'h1112: d <= 8'hC0; 15'h1113: d <= 8'hC0;
                15'h1114: d <= 8'hC0; 15'h1115: d <= 8'hC0; 15'h1116: d <= 8'hC0; 15'h1117: d <= 8'hC0;
                15'h1118: d <= 8'hC0; 15'h1119: d <= 8'hC0; 15'h111A: d <= 8'hC0; 15'h111B: d <= 8'hC0;
                15'h111C: d <= 8'hC0; 15'h111D: d <= 8'hC0; 15'h111E: d <= 8'hC0; 15'h111F: d <= 8'hC0;
                15'h1120: d <= 8'hC0; 15'h1121: d <= 8'hC0; 15'h1122: d <= 8'hC0; 15'h1123: d <= 8'hC0;
                15'h1124: d <= 8'hC0; 15'h1125: d <= 8'hC0; 15'h1126: d <= 8'hC0; 15'h1127: d <= 8'hC0;
                15'h1128: d <= 8'hC0; 15'h1129: d <= 8'hC0; 15'h112A: d <= 8'hC0; 15'h112B: d <= 8'hC0;
                15'h112C: d <= 8'hC0; 15'h112D: d <= 8'hC0; 15'h112E: d <= 8'hC0; 15'h112F: d <= 8'hC0;
                15'h1130: d <= 8'hC0; 15'h1131: d <= 8'hC0; 15'h1132: d <= 8'hC0; 15'h1133: d <= 8'hC0;
                15'h1134: d <= 8'hC0; 15'h1135: d <= 8'hC0; 15'h1136: d <= 8'hC0; 15'h1137: d <= 8'hC0;
                15'h1138: d <= 8'hC0; 15'h1139: d <= 8'hC0; 15'h113A: d <= 8'hC0; 15'h113B: d <= 8'hC0;
                15'h113C: d <= 8'hC0; 15'h113D: d <= 8'hC0; 15'h113E: d <= 8'hC0; 15'h113F: d <= 8'hC0;
                15'h1140: d <= 8'hC0; 15'h1141: d <= 8'hC0; 15'h1142: d <= 8'hC0; 15'h1143: d <= 8'hC0;
                15'h1144: d <= 8'hC0; 15'h1145: d <= 8'hC0; 15'h1146: d <= 8'hC0; 15'h1147: d <= 8'hC0;
                15'h1148: d <= 8'hC0; 15'h1149: d <= 8'hC0; 15'h114A: d <= 8'hC0; 15'h114B: d <= 8'hC0;
                15'h114C: d <= 8'hC0; 15'h114D: d <= 8'hC0; 15'h114E: d <= 8'hC0; 15'h114F: d <= 8'hC0;
                15'h1150: d <= 8'hC0; 15'h1151: d <= 8'hC0; 15'h1152: d <= 8'hC0; 15'h1153: d <= 8'hC0;
                15'h1154: d <= 8'hC0; 15'h1155: d <= 8'hC0; 15'h1156: d <= 8'hC0; 15'h1157: d <= 8'hC0;
                15'h1158: d <= 8'hC0; 15'h1159: d <= 8'hC0; 15'h115A: d <= 8'hC0; 15'h115B: d <= 8'hC0;
                15'h115C: d <= 8'hC0; 15'h115D: d <= 8'hC0; 15'h115E: d <= 8'hC0; 15'h115F: d <= 8'hC0;
                15'h1160: d <= 8'hC0; 15'h1161: d <= 8'hC0; 15'h1162: d <= 8'hC0; 15'h1163: d <= 8'hC0;
                15'h1164: d <= 8'hC0; 15'h1165: d <= 8'hC0; 15'h1166: d <= 8'hC0; 15'h1167: d <= 8'hC0;
                15'h1168: d <= 8'hC0; 15'h1169: d <= 8'hC0; 15'h116A: d <= 8'hC0; 15'h116B: d <= 8'hC0;
                15'h116C: d <= 8'hC0; 15'h116D: d <= 8'hC0; 15'h116E: d <= 8'hC0; 15'h116F: d <= 8'hC0;
                15'h1170: d <= 8'hC0; 15'h1171: d <= 8'hC0; 15'h1172: d <= 8'hC0; 15'h1173: d <= 8'hC0;
                15'h1174: d <= 8'hC0; 15'h1175: d <= 8'hC0; 15'h1176: d <= 8'hC0; 15'h1177: d <= 8'hC0;
                15'h1178: d <= 8'hC0; 15'h1179: d <= 8'hC0; 15'h117A: d <= 8'hC0; 15'h117B: d <= 8'hC0;
                15'h117C: d <= 8'hC0; 15'h117D: d <= 8'hC0; 15'h117E: d <= 8'hC0; 15'h117F: d <= 8'hC0;
                15'h1180: d <= 8'hC0; 15'h1181: d <= 8'hC0; 15'h1182: d <= 8'hC0; 15'h1183: d <= 8'hC0;
                15'h1184: d <= 8'hC0; 15'h1185: d <= 8'hC0; 15'h1186: d <= 8'hC0; 15'h1187: d <= 8'hC0;
                15'h1188: d <= 8'hC0; 15'h1189: d <= 8'hC0; 15'h118A: d <= 8'hC0; 15'h118B: d <= 8'hC0;
                15'h118C: d <= 8'hC0; 15'h118D: d <= 8'hC0; 15'h118E: d <= 8'hC0; 15'h118F: d <= 8'hC0;
                15'h1190: d <= 8'hC0; 15'h1191: d <= 8'hC0; 15'h1192: d <= 8'hC0; 15'h1193: d <= 8'hC0;
                15'h1194: d <= 8'hC0; 15'h1195: d <= 8'hC0; 15'h1196: d <= 8'hC0; 15'h1197: d <= 8'hC0;
                15'h1198: d <= 8'hC0; 15'h1199: d <= 8'hC0; 15'h119A: d <= 8'hC0; 15'h119B: d <= 8'hC0;
                15'h119C: d <= 8'hC0; 15'h119D: d <= 8'hC0; 15'h119E: d <= 8'hC0; 15'h119F: d <= 8'hC0;
                15'h11A0: d <= 8'hC0; 15'h11A1: d <= 8'hC0; 15'h11A2: d <= 8'hC0; 15'h11A3: d <= 8'hC0;
                15'h11A4: d <= 8'hC0; 15'h11A5: d <= 8'hC0; 15'h11A6: d <= 8'hC0; 15'h11A7: d <= 8'hC0;
                15'h11A8: d <= 8'hC0; 15'h11A9: d <= 8'hC0; 15'h11AA: d <= 8'hC0; 15'h11AB: d <= 8'hC0;
                15'h11AC: d <= 8'hC0; 15'h11AD: d <= 8'hC0; 15'h11AE: d <= 8'hC0; 15'h11AF: d <= 8'hC0;
                15'h11B0: d <= 8'hC0; 15'h11B1: d <= 8'hC0; 15'h11B2: d <= 8'hC0; 15'h11B3: d <= 8'hC0;
                15'h11B4: d <= 8'hC0; 15'h11B5: d <= 8'hC0; 15'h11B6: d <= 8'hC0; 15'h11B7: d <= 8'hC0;
                15'h11B8: d <= 8'hC0; 15'h11B9: d <= 8'hC0; 15'h11BA: d <= 8'hC0; 15'h11BB: d <= 8'hC0;
                15'h11BC: d <= 8'hC0; 15'h11BD: d <= 8'hC0; 15'h11BE: d <= 8'hC0; 15'h11BF: d <= 8'hC0;
                15'h11C0: d <= 8'hC0; 15'h11C1: d <= 8'hC0; 15'h11C2: d <= 8'hC0; 15'h11C3: d <= 8'hC0;
                15'h11C4: d <= 8'hC0; 15'h11C5: d <= 8'hC0; 15'h11C6: d <= 8'hC0; 15'h11C7: d <= 8'hC0;
                15'h11C8: d <= 8'hC0; 15'h11C9: d <= 8'hC0; 15'h11CA: d <= 8'hC0; 15'h11CB: d <= 8'hC0;
                15'h11CC: d <= 8'hC0; 15'h11CD: d <= 8'hC0; 15'h11CE: d <= 8'hC0; 15'h11CF: d <= 8'hC0;
                15'h11D0: d <= 8'hC0; 15'h11D1: d <= 8'hC0; 15'h11D2: d <= 8'hC0; 15'h11D3: d <= 8'hC0;
                15'h11D4: d <= 8'hC0; 15'h11D5: d <= 8'hC0; 15'h11D6: d <= 8'hC0; 15'h11D7: d <= 8'hC0;
                15'h11D8: d <= 8'hC0; 15'h11D9: d <= 8'hC0; 15'h11DA: d <= 8'hC0; 15'h11DB: d <= 8'hC0;
                15'h11DC: d <= 8'hC0; 15'h11DD: d <= 8'hC0; 15'h11DE: d <= 8'hC0; 15'h11DF: d <= 8'hC0;
                15'h11E0: d <= 8'hC0; 15'h11E1: d <= 8'hC0; 15'h11E2: d <= 8'hC0; 15'h11E3: d <= 8'hC0;
                15'h11E4: d <= 8'hC0; 15'h11E5: d <= 8'hC0; 15'h11E6: d <= 8'hC0; 15'h11E7: d <= 8'hC0;
                15'h11E8: d <= 8'hC0; 15'h11E9: d <= 8'hC0; 15'h11EA: d <= 8'hC0; 15'h11EB: d <= 8'hC0;
                15'h11EC: d <= 8'hC0; 15'h11ED: d <= 8'hC0; 15'h11EE: d <= 8'hC0; 15'h11EF: d <= 8'hC0;
                15'h11F0: d <= 8'hC0; 15'h11F1: d <= 8'hC0; 15'h11F2: d <= 8'hC0; 15'h11F3: d <= 8'hC0;
                15'h11F4: d <= 8'hC0; 15'h11F5: d <= 8'hC0; 15'h11F6: d <= 8'hC0; 15'h11F7: d <= 8'hC0;
                15'h11F8: d <= 8'hC0; 15'h11F9: d <= 8'hC0; 15'h11FA: d <= 8'hC0; 15'h11FB: d <= 8'hC0;
                15'h11FC: d <= 8'hC0; 15'h11FD: d <= 8'hC0; 15'h11FE: d <= 8'hC0; 15'h11FF: d <= 8'hC0;
                15'h1200: d <= 8'hC0; 15'h1201: d <= 8'hC0; 15'h1202: d <= 8'hC0; 15'h1203: d <= 8'hC0;
                15'h1204: d <= 8'hC0; 15'h1205: d <= 8'hC0; 15'h1206: d <= 8'hC0; 15'h1207: d <= 8'hC0;
                15'h1208: d <= 8'hC0; 15'h1209: d <= 8'hC0; 15'h120A: d <= 8'hC0; 15'h120B: d <= 8'hC0;
                15'h120C: d <= 8'hC0; 15'h120D: d <= 8'hC0; 15'h120E: d <= 8'hC0; 15'h120F: d <= 8'hC0;
                15'h1210: d <= 8'hC0; 15'h1211: d <= 8'hC0; 15'h1212: d <= 8'hC0; 15'h1213: d <= 8'hC0;
                15'h1214: d <= 8'hC0; 15'h1215: d <= 8'hC0; 15'h1216: d <= 8'hC0; 15'h1217: d <= 8'hC0;
                15'h1218: d <= 8'hC0; 15'h1219: d <= 8'hC0; 15'h121A: d <= 8'hC0; 15'h121B: d <= 8'hC0;
                15'h121C: d <= 8'hC0; 15'h121D: d <= 8'hC0; 15'h121E: d <= 8'hC0; 15'h121F: d <= 8'hC0;
                15'h1220: d <= 8'hC0; 15'h1221: d <= 8'hC0; 15'h1222: d <= 8'hC0; 15'h1223: d <= 8'hC0;
                15'h1224: d <= 8'hC0; 15'h1225: d <= 8'hC0; 15'h1226: d <= 8'hC0; 15'h1227: d <= 8'hC0;
                15'h1228: d <= 8'hC0; 15'h1229: d <= 8'hC0; 15'h122A: d <= 8'hC0; 15'h122B: d <= 8'hC0;
                15'h122C: d <= 8'hC0; 15'h122D: d <= 8'hC0; 15'h122E: d <= 8'hC0; 15'h122F: d <= 8'hC0;
                15'h1230: d <= 8'hC0; 15'h1231: d <= 8'hC0; 15'h1232: d <= 8'hC0; 15'h1233: d <= 8'hC0;
                15'h1234: d <= 8'hC0; 15'h1235: d <= 8'hC0; 15'h1236: d <= 8'hC0; 15'h1237: d <= 8'hC0;
                15'h1238: d <= 8'hC0; 15'h1239: d <= 8'hC0; 15'h123A: d <= 8'hC0; 15'h123B: d <= 8'hC0;
                15'h123C: d <= 8'hC0; 15'h123D: d <= 8'hC0; 15'h123E: d <= 8'hC0; 15'h123F: d <= 8'hC0;
                15'h1240: d <= 8'hC0; 15'h1241: d <= 8'hC0; 15'h1242: d <= 8'hC0; 15'h1243: d <= 8'hC0;
                15'h1244: d <= 8'hC0; 15'h1245: d <= 8'hC0; 15'h1246: d <= 8'hC0; 15'h1247: d <= 8'hC0;
                15'h1248: d <= 8'hC0; 15'h1249: d <= 8'hC0; 15'h124A: d <= 8'hC0; 15'h124B: d <= 8'hC0;
                15'h124C: d <= 8'hC0; 15'h124D: d <= 8'hC0; 15'h124E: d <= 8'hC0; 15'h124F: d <= 8'hC0;
                15'h1250: d <= 8'hC0; 15'h1251: d <= 8'hC0; 15'h1252: d <= 8'hC0; 15'h1253: d <= 8'hC0;
                15'h1254: d <= 8'hC0; 15'h1255: d <= 8'hC0; 15'h1256: d <= 8'hC0; 15'h1257: d <= 8'hC0;
                15'h1258: d <= 8'hC0; 15'h1259: d <= 8'hC0; 15'h125A: d <= 8'hC0; 15'h125B: d <= 8'hC0;
                15'h125C: d <= 8'hC0; 15'h125D: d <= 8'hC0; 15'h125E: d <= 8'hC0; 15'h125F: d <= 8'hC0;
                15'h1260: d <= 8'hC0; 15'h1261: d <= 8'hC0; 15'h1262: d <= 8'hC0; 15'h1263: d <= 8'hC0;
                15'h1264: d <= 8'hC0; 15'h1265: d <= 8'hC0; 15'h1266: d <= 8'hC0; 15'h1267: d <= 8'hC0;
                15'h1268: d <= 8'hC0; 15'h1269: d <= 8'hC0; 15'h126A: d <= 8'hC0; 15'h126B: d <= 8'hC0;
                15'h126C: d <= 8'hC0; 15'h126D: d <= 8'hC0; 15'h126E: d <= 8'hC0; 15'h126F: d <= 8'hC0;
                15'h1270: d <= 8'hC0; 15'h1271: d <= 8'hC0; 15'h1272: d <= 8'hC0; 15'h1273: d <= 8'hC0;
                15'h1274: d <= 8'hC0; 15'h1275: d <= 8'hC0; 15'h1276: d <= 8'hC0; 15'h1277: d <= 8'hC0;
                15'h1278: d <= 8'hC0; 15'h1279: d <= 8'hC0; 15'h127A: d <= 8'hC0; 15'h127B: d <= 8'hC0;
                15'h127C: d <= 8'hC0; 15'h127D: d <= 8'hC0; 15'h127E: d <= 8'hC0; 15'h127F: d <= 8'hC0;
                15'h1280: d <= 8'hC0; 15'h1281: d <= 8'hC0; 15'h1282: d <= 8'hC0; 15'h1283: d <= 8'hC0;
                15'h1284: d <= 8'hC0; 15'h1285: d <= 8'hC0; 15'h1286: d <= 8'hC0; 15'h1287: d <= 8'hC0;
                15'h1288: d <= 8'hC0; 15'h1289: d <= 8'hC0; 15'h128A: d <= 8'hC0; 15'h128B: d <= 8'hC0;
                15'h128C: d <= 8'hC0; 15'h128D: d <= 8'hC0; 15'h128E: d <= 8'hC0; 15'h128F: d <= 8'hC0;
                15'h1290: d <= 8'hC0; 15'h1291: d <= 8'hC0; 15'h1292: d <= 8'hC0; 15'h1293: d <= 8'hC0;
                15'h1294: d <= 8'hC0; 15'h1295: d <= 8'hC0; 15'h1296: d <= 8'hC0; 15'h1297: d <= 8'hC0;
                15'h1298: d <= 8'hC0; 15'h1299: d <= 8'hC0; 15'h129A: d <= 8'hC0; 15'h129B: d <= 8'hC0;
                15'h129C: d <= 8'hC0; 15'h129D: d <= 8'hC0; 15'h129E: d <= 8'hC0; 15'h129F: d <= 8'hC0;
                15'h12A0: d <= 8'hC0; 15'h12A1: d <= 8'hC0; 15'h12A2: d <= 8'hC0; 15'h12A3: d <= 8'hC0;
                15'h12A4: d <= 8'hC0; 15'h12A5: d <= 8'hC0; 15'h12A6: d <= 8'hC0; 15'h12A7: d <= 8'hC0;
                15'h12A8: d <= 8'hC0; 15'h12A9: d <= 8'hC0; 15'h12AA: d <= 8'hC0; 15'h12AB: d <= 8'hC0;
                15'h12AC: d <= 8'hC0; 15'h12AD: d <= 8'hC0; 15'h12AE: d <= 8'hC0; 15'h12AF: d <= 8'hC0;
                15'h12B0: d <= 8'hC0; 15'h12B1: d <= 8'hC0; 15'h12B2: d <= 8'hC0; 15'h12B3: d <= 8'hC0;
                15'h12B4: d <= 8'hC0; 15'h12B5: d <= 8'hC0; 15'h12B6: d <= 8'hC0; 15'h12B7: d <= 8'hC0;
                15'h12B8: d <= 8'hC0; 15'h12B9: d <= 8'hC0; 15'h12BA: d <= 8'hC0; 15'h12BB: d <= 8'hC0;
                15'h12BC: d <= 8'hC0; 15'h12BD: d <= 8'hC0; 15'h12BE: d <= 8'hC0; 15'h12BF: d <= 8'hC0;
                15'h12C0: d <= 8'hC0; 15'h12C1: d <= 8'hC0; 15'h12C2: d <= 8'hC0; 15'h12C3: d <= 8'hC0;
                15'h12C4: d <= 8'hC0; 15'h12C5: d <= 8'hC0; 15'h12C6: d <= 8'hC0; 15'h12C7: d <= 8'hC0;
                15'h12C8: d <= 8'hC0; 15'h12C9: d <= 8'hC0; 15'h12CA: d <= 8'hC0; 15'h12CB: d <= 8'hC0;
                15'h12CC: d <= 8'hC0; 15'h12CD: d <= 8'hC0; 15'h12CE: d <= 8'hC0; 15'h12CF: d <= 8'hC0;
                15'h12D0: d <= 8'hC0; 15'h12D1: d <= 8'hC0; 15'h12D2: d <= 8'hC0; 15'h12D3: d <= 8'hC0;
                15'h12D4: d <= 8'hC0; 15'h12D5: d <= 8'hC0; 15'h12D6: d <= 8'hC0; 15'h12D7: d <= 8'hC0;
                15'h12D8: d <= 8'hC0; 15'h12D9: d <= 8'hC0; 15'h12DA: d <= 8'hC0; 15'h12DB: d <= 8'hC0;
                15'h12DC: d <= 8'hC0; 15'h12DD: d <= 8'hC0; 15'h12DE: d <= 8'hC0; 15'h12DF: d <= 8'hC0;
                15'h12E0: d <= 8'hC0; 15'h12E1: d <= 8'hC0; 15'h12E2: d <= 8'hC0; 15'h12E3: d <= 8'hC0;
                15'h12E4: d <= 8'hC0; 15'h12E5: d <= 8'hC0; 15'h12E6: d <= 8'hC0; 15'h12E7: d <= 8'hC0;
                15'h12E8: d <= 8'hC0; 15'h12E9: d <= 8'hC0; 15'h12EA: d <= 8'hC0; 15'h12EB: d <= 8'hC0;
                15'h12EC: d <= 8'hC0; 15'h12ED: d <= 8'hC0; 15'h12EE: d <= 8'hC0; 15'h12EF: d <= 8'hC0;
                15'h12F0: d <= 8'hC0; 15'h12F1: d <= 8'hC0; 15'h12F2: d <= 8'hC0; 15'h12F3: d <= 8'hC0;
                15'h12F4: d <= 8'hC0; 15'h12F5: d <= 8'hC0; 15'h12F6: d <= 8'hC0; 15'h12F7: d <= 8'hC0;
                15'h12F8: d <= 8'hC0; 15'h12F9: d <= 8'hC0; 15'h12FA: d <= 8'hC0; 15'h12FB: d <= 8'hC0;
                15'h12FC: d <= 8'hC0; 15'h12FD: d <= 8'hC0; 15'h12FE: d <= 8'hC0; 15'h12FF: d <= 8'hC0;
                15'h1300: d <= 8'hC0; 15'h1301: d <= 8'hC0; 15'h1302: d <= 8'hC0; 15'h1303: d <= 8'hC0;
                15'h1304: d <= 8'hC0; 15'h1305: d <= 8'hC0; 15'h1306: d <= 8'hC0; 15'h1307: d <= 8'hC0;
                15'h1308: d <= 8'hC0; 15'h1309: d <= 8'hC0; 15'h130A: d <= 8'hC0; 15'h130B: d <= 8'hC0;
                15'h130C: d <= 8'hC0; 15'h130D: d <= 8'hC0; 15'h130E: d <= 8'hC0; 15'h130F: d <= 8'hC0;
                15'h1310: d <= 8'hC0; 15'h1311: d <= 8'hC0; 15'h1312: d <= 8'hC0; 15'h1313: d <= 8'hC0;
                15'h1314: d <= 8'hC0; 15'h1315: d <= 8'hC0; 15'h1316: d <= 8'hC0; 15'h1317: d <= 8'hC0;
                15'h1318: d <= 8'hC0; 15'h1319: d <= 8'hC0; 15'h131A: d <= 8'hC0; 15'h131B: d <= 8'hC0;
                15'h131C: d <= 8'hC0; 15'h131D: d <= 8'hC0; 15'h131E: d <= 8'hC0; 15'h131F: d <= 8'hC0;
                15'h1320: d <= 8'hC0; 15'h1321: d <= 8'hC0; 15'h1322: d <= 8'hC0; 15'h1323: d <= 8'hC0;
                15'h1324: d <= 8'hC0; 15'h1325: d <= 8'hC0; 15'h1326: d <= 8'hC0; 15'h1327: d <= 8'hC0;
                15'h1328: d <= 8'hC0; 15'h1329: d <= 8'hC0; 15'h132A: d <= 8'hC0; 15'h132B: d <= 8'hC0;
                15'h132C: d <= 8'hC0; 15'h132D: d <= 8'hC0; 15'h132E: d <= 8'hC0; 15'h132F: d <= 8'hC0;
                15'h1330: d <= 8'hC0; 15'h1331: d <= 8'hC0; 15'h1332: d <= 8'hC0; 15'h1333: d <= 8'hC0;
                15'h1334: d <= 8'hC0; 15'h1335: d <= 8'hC0; 15'h1336: d <= 8'hC0; 15'h1337: d <= 8'hC0;
                15'h1338: d <= 8'hC0; 15'h1339: d <= 8'hC0; 15'h133A: d <= 8'hC0; 15'h133B: d <= 8'hC0;
                15'h133C: d <= 8'hC0; 15'h133D: d <= 8'hC0; 15'h133E: d <= 8'hC0; 15'h133F: d <= 8'hC0;
                15'h1340: d <= 8'hC0; 15'h1341: d <= 8'hC0; 15'h1342: d <= 8'hC0; 15'h1343: d <= 8'hC0;
                15'h1344: d <= 8'hC0; 15'h1345: d <= 8'hC0; 15'h1346: d <= 8'hC0; 15'h1347: d <= 8'hC0;
                15'h1348: d <= 8'hC0; 15'h1349: d <= 8'hC0; 15'h134A: d <= 8'hC0; 15'h134B: d <= 8'hC0;
                15'h134C: d <= 8'hC0; 15'h134D: d <= 8'hC0; 15'h134E: d <= 8'hC0; 15'h134F: d <= 8'hC0;
                15'h1350: d <= 8'hC0; 15'h1351: d <= 8'hC0; 15'h1352: d <= 8'hC0; 15'h1353: d <= 8'hC0;
                15'h1354: d <= 8'hC0; 15'h1355: d <= 8'hC0; 15'h1356: d <= 8'hC0; 15'h1357: d <= 8'hC0;
                15'h1358: d <= 8'hC0; 15'h1359: d <= 8'hC0; 15'h135A: d <= 8'hC0; 15'h135B: d <= 8'hC0;
                15'h135C: d <= 8'hC0; 15'h135D: d <= 8'hC0; 15'h135E: d <= 8'hC0; 15'h135F: d <= 8'hC0;
                15'h1360: d <= 8'hC0; 15'h1361: d <= 8'hC0; 15'h1362: d <= 8'hC0; 15'h1363: d <= 8'hC0;
                15'h1364: d <= 8'hC0; 15'h1365: d <= 8'hC0; 15'h1366: d <= 8'hC0; 15'h1367: d <= 8'hC0;
                15'h1368: d <= 8'hC0; 15'h1369: d <= 8'hC0; 15'h136A: d <= 8'hC0; 15'h136B: d <= 8'hC0;
                15'h136C: d <= 8'hC0; 15'h136D: d <= 8'hC0; 15'h136E: d <= 8'hC0; 15'h136F: d <= 8'hC0;
                15'h1370: d <= 8'hC0; 15'h1371: d <= 8'hC0; 15'h1372: d <= 8'hC0; 15'h1373: d <= 8'hC0;
                15'h1374: d <= 8'hC0; 15'h1375: d <= 8'hC0; 15'h1376: d <= 8'hC0; 15'h1377: d <= 8'hC0;
                15'h1378: d <= 8'hC0; 15'h1379: d <= 8'hC0; 15'h137A: d <= 8'hC0; 15'h137B: d <= 8'hC0;
                15'h137C: d <= 8'hC0; 15'h137D: d <= 8'hC0; 15'h137E: d <= 8'hC0; 15'h137F: d <= 8'hC0;
                15'h1380: d <= 8'hC0; 15'h1381: d <= 8'hC0; 15'h1382: d <= 8'hC0; 15'h1383: d <= 8'hC0;
                15'h1384: d <= 8'hC0; 15'h1385: d <= 8'hC0; 15'h1386: d <= 8'hC0; 15'h1387: d <= 8'hC0;
                15'h1388: d <= 8'hC0; 15'h1389: d <= 8'hC0; 15'h138A: d <= 8'hC0; 15'h138B: d <= 8'hC0;
                15'h138C: d <= 8'hC0; 15'h138D: d <= 8'hC0; 15'h138E: d <= 8'hC0; 15'h138F: d <= 8'hC0;
                15'h1390: d <= 8'hC0; 15'h1391: d <= 8'hC0; 15'h1392: d <= 8'hC0; 15'h1393: d <= 8'hC0;
                15'h1394: d <= 8'hC0; 15'h1395: d <= 8'hC0; 15'h1396: d <= 8'hC0; 15'h1397: d <= 8'hC0;
                15'h1398: d <= 8'hC0; 15'h1399: d <= 8'hC0; 15'h139A: d <= 8'hC0; 15'h139B: d <= 8'hC0;
                15'h139C: d <= 8'hC0; 15'h139D: d <= 8'hC0; 15'h139E: d <= 8'hC0; 15'h139F: d <= 8'hC0;
                15'h13A0: d <= 8'hC0; 15'h13A1: d <= 8'hC0; 15'h13A2: d <= 8'hC0; 15'h13A3: d <= 8'hC0;
                15'h13A4: d <= 8'hC0; 15'h13A5: d <= 8'hC0; 15'h13A6: d <= 8'hC0; 15'h13A7: d <= 8'hC0;
                15'h13A8: d <= 8'hC0; 15'h13A9: d <= 8'hC0; 15'h13AA: d <= 8'hC0; 15'h13AB: d <= 8'hC0;
                15'h13AC: d <= 8'hC0; 15'h13AD: d <= 8'hC0; 15'h13AE: d <= 8'hC0; 15'h13AF: d <= 8'hC0;
                15'h13B0: d <= 8'hC0; 15'h13B1: d <= 8'hC0; 15'h13B2: d <= 8'hC0; 15'h13B3: d <= 8'hC0;
                15'h13B4: d <= 8'hC0; 15'h13B5: d <= 8'hC0; 15'h13B6: d <= 8'hC0; 15'h13B7: d <= 8'hC0;
                15'h13B8: d <= 8'hC0; 15'h13B9: d <= 8'hC0; 15'h13BA: d <= 8'hC0; 15'h13BB: d <= 8'hC0;
                15'h13BC: d <= 8'hC0; 15'h13BD: d <= 8'hC0; 15'h13BE: d <= 8'hC0; 15'h13BF: d <= 8'hC0;
                15'h13C0: d <= 8'hC0; 15'h13C1: d <= 8'hC0; 15'h13C2: d <= 8'hC0; 15'h13C3: d <= 8'hC0;
                15'h13C4: d <= 8'hC0; 15'h13C5: d <= 8'hC0; 15'h13C6: d <= 8'hC0; 15'h13C7: d <= 8'hC0;
                15'h13C8: d <= 8'hC0; 15'h13C9: d <= 8'hC0; 15'h13CA: d <= 8'hC0; 15'h13CB: d <= 8'hC0;
                15'h13CC: d <= 8'hC0; 15'h13CD: d <= 8'hC0; 15'h13CE: d <= 8'hC0; 15'h13CF: d <= 8'hC0;
                15'h13D0: d <= 8'hC0; 15'h13D1: d <= 8'hC0; 15'h13D2: d <= 8'hC0; 15'h13D3: d <= 8'hC0;
                15'h13D4: d <= 8'hC0; 15'h13D5: d <= 8'hC0; 15'h13D6: d <= 8'hC0; 15'h13D7: d <= 8'hC0;
                15'h13D8: d <= 8'hC0; 15'h13D9: d <= 8'hC0; 15'h13DA: d <= 8'hC0; 15'h13DB: d <= 8'hC0;
                15'h13DC: d <= 8'hC0; 15'h13DD: d <= 8'hC0; 15'h13DE: d <= 8'hC0; 15'h13DF: d <= 8'hC0;
                15'h13E0: d <= 8'hC0; 15'h13E1: d <= 8'hC0; 15'h13E2: d <= 8'hC0; 15'h13E3: d <= 8'hC0;
                15'h13E4: d <= 8'hC0; 15'h13E5: d <= 8'hC0; 15'h13E6: d <= 8'hC0; 15'h13E7: d <= 8'hC0;
                15'h13E8: d <= 8'hC0; 15'h13E9: d <= 8'hC0; 15'h13EA: d <= 8'hC0; 15'h13EB: d <= 8'hC0;
                15'h13EC: d <= 8'hC0; 15'h13ED: d <= 8'hC0; 15'h13EE: d <= 8'hC0; 15'h13EF: d <= 8'hC0;
                15'h13F0: d <= 8'hC0; 15'h13F1: d <= 8'hC0; 15'h13F2: d <= 8'hC0; 15'h13F3: d <= 8'hC0;
                15'h13F4: d <= 8'hC0; 15'h13F5: d <= 8'hC0; 15'h13F6: d <= 8'hC0; 15'h13F7: d <= 8'hC0;
                15'h13F8: d <= 8'hC0; 15'h13F9: d <= 8'hC0; 15'h13FA: d <= 8'hC0; 15'h13FB: d <= 8'hC0;
                15'h13FC: d <= 8'hC0; 15'h13FD: d <= 8'hC0; 15'h13FE: d <= 8'hC0; 15'h13FF: d <= 8'hC0;
                15'h1400: d <= 8'hC0; 15'h1401: d <= 8'hC0; 15'h1402: d <= 8'hC0; 15'h1403: d <= 8'hC0;
                15'h1404: d <= 8'hC0; 15'h1405: d <= 8'hC0; 15'h1406: d <= 8'hC0; 15'h1407: d <= 8'hC0;
                15'h1408: d <= 8'hC0; 15'h1409: d <= 8'hC0; 15'h140A: d <= 8'hC0; 15'h140B: d <= 8'hC0;
                15'h140C: d <= 8'hC0; 15'h140D: d <= 8'hC0; 15'h140E: d <= 8'hC0; 15'h140F: d <= 8'hC0;
                15'h1410: d <= 8'hC0; 15'h1411: d <= 8'hC0; 15'h1412: d <= 8'hC0; 15'h1413: d <= 8'hC0;
                15'h1414: d <= 8'hC0; 15'h1415: d <= 8'hC0; 15'h1416: d <= 8'hC0; 15'h1417: d <= 8'hC0;
                15'h1418: d <= 8'hC0; 15'h1419: d <= 8'hC0; 15'h141A: d <= 8'hC0; 15'h141B: d <= 8'hC0;
                15'h141C: d <= 8'hC0; 15'h141D: d <= 8'hC0; 15'h141E: d <= 8'hC0; 15'h141F: d <= 8'hC0;
                15'h1420: d <= 8'hC0; 15'h1421: d <= 8'hC0; 15'h1422: d <= 8'hC0; 15'h1423: d <= 8'hC0;
                15'h1424: d <= 8'hC0; 15'h1425: d <= 8'hC0; 15'h1426: d <= 8'hC0; 15'h1427: d <= 8'hC0;
                15'h1428: d <= 8'hC0; 15'h1429: d <= 8'hC0; 15'h142A: d <= 8'hC0; 15'h142B: d <= 8'hC0;
                15'h142C: d <= 8'hC0; 15'h142D: d <= 8'hC0; 15'h142E: d <= 8'hC0; 15'h142F: d <= 8'hC0;
                15'h1430: d <= 8'hC0; 15'h1431: d <= 8'hC0; 15'h1432: d <= 8'hC0; 15'h1433: d <= 8'hC0;
                15'h1434: d <= 8'hC0; 15'h1435: d <= 8'hC0; 15'h1436: d <= 8'hC0; 15'h1437: d <= 8'hC0;
                15'h1438: d <= 8'hC0; 15'h1439: d <= 8'hC0; 15'h143A: d <= 8'hC0; 15'h143B: d <= 8'hC0;
                15'h143C: d <= 8'hC0; 15'h143D: d <= 8'hC0; 15'h143E: d <= 8'hC0; 15'h143F: d <= 8'hC0;
                15'h1440: d <= 8'hC0; 15'h1441: d <= 8'hC0; 15'h1442: d <= 8'hC0; 15'h1443: d <= 8'hC0;
                15'h1444: d <= 8'hC0; 15'h1445: d <= 8'hC0; 15'h1446: d <= 8'hC0; 15'h1447: d <= 8'hC0;
                15'h1448: d <= 8'hC0; 15'h1449: d <= 8'hC0; 15'h144A: d <= 8'hC0; 15'h144B: d <= 8'hC0;
                15'h144C: d <= 8'hC0; 15'h144D: d <= 8'hC0; 15'h144E: d <= 8'hC0; 15'h144F: d <= 8'hC0;
                15'h1450: d <= 8'hC0; 15'h1451: d <= 8'hC0; 15'h1452: d <= 8'hC0; 15'h1453: d <= 8'hC0;
                15'h1454: d <= 8'hC0; 15'h1455: d <= 8'hC0; 15'h1456: d <= 8'hC0; 15'h1457: d <= 8'hC0;
                15'h1458: d <= 8'hC0; 15'h1459: d <= 8'hC0; 15'h145A: d <= 8'hC0; 15'h145B: d <= 8'hC0;
                15'h145C: d <= 8'hC0; 15'h145D: d <= 8'hC0; 15'h145E: d <= 8'hC0; 15'h145F: d <= 8'hC0;
                15'h1460: d <= 8'hC0; 15'h1461: d <= 8'hC0; 15'h1462: d <= 8'hC0; 15'h1463: d <= 8'hC0;
                15'h1464: d <= 8'hC0; 15'h1465: d <= 8'hC0; 15'h1466: d <= 8'hC0; 15'h1467: d <= 8'hC0;
                15'h1468: d <= 8'hC0; 15'h1469: d <= 8'hC0; 15'h146A: d <= 8'hC0; 15'h146B: d <= 8'hC0;
                15'h146C: d <= 8'hC0; 15'h146D: d <= 8'hC0; 15'h146E: d <= 8'hC0; 15'h146F: d <= 8'hC0;
                15'h1470: d <= 8'hC0; 15'h1471: d <= 8'hC0; 15'h1472: d <= 8'hC0; 15'h1473: d <= 8'hC0;
                15'h1474: d <= 8'hC0; 15'h1475: d <= 8'hC0; 15'h1476: d <= 8'hC0; 15'h1477: d <= 8'hC0;
                15'h1478: d <= 8'hC0; 15'h1479: d <= 8'hC0; 15'h147A: d <= 8'hC0; 15'h147B: d <= 8'hC0;
                15'h147C: d <= 8'hC0; 15'h147D: d <= 8'hC0; 15'h147E: d <= 8'hC0; 15'h147F: d <= 8'hC0;
                15'h1480: d <= 8'hC0; 15'h1481: d <= 8'hC0; 15'h1482: d <= 8'hC0; 15'h1483: d <= 8'hC0;
                15'h1484: d <= 8'hC0; 15'h1485: d <= 8'hC0; 15'h1486: d <= 8'hC0; 15'h1487: d <= 8'hC0;
                15'h1488: d <= 8'hC0; 15'h1489: d <= 8'hC0; 15'h148A: d <= 8'hC0; 15'h148B: d <= 8'hC0;
                15'h148C: d <= 8'hC0; 15'h148D: d <= 8'hC0; 15'h148E: d <= 8'hC0; 15'h148F: d <= 8'hC0;
                15'h1490: d <= 8'hC0; 15'h1491: d <= 8'hC0; 15'h1492: d <= 8'hC0; 15'h1493: d <= 8'hC0;
                15'h1494: d <= 8'hC0; 15'h1495: d <= 8'hC0; 15'h1496: d <= 8'hC0; 15'h1497: d <= 8'hC0;
                15'h1498: d <= 8'hC0; 15'h1499: d <= 8'hC0; 15'h149A: d <= 8'hC0; 15'h149B: d <= 8'hC0;
                15'h149C: d <= 8'hC0; 15'h149D: d <= 8'hC0; 15'h149E: d <= 8'hC0; 15'h149F: d <= 8'hC0;
                15'h14A0: d <= 8'hC0; 15'h14A1: d <= 8'hC0; 15'h14A2: d <= 8'hC0; 15'h14A3: d <= 8'hC0;
                15'h14A4: d <= 8'hC0; 15'h14A5: d <= 8'hC0; 15'h14A6: d <= 8'hC0; 15'h14A7: d <= 8'hC0;
                15'h14A8: d <= 8'hC0; 15'h14A9: d <= 8'hC0; 15'h14AA: d <= 8'hC0; 15'h14AB: d <= 8'hC0;
                15'h14AC: d <= 8'hC0; 15'h14AD: d <= 8'hC0; 15'h14AE: d <= 8'hC0; 15'h14AF: d <= 8'hC0;
                15'h14B0: d <= 8'hC0; 15'h14B1: d <= 8'hC0; 15'h14B2: d <= 8'hC0; 15'h14B3: d <= 8'hC0;
                15'h14B4: d <= 8'hC0; 15'h14B5: d <= 8'hC0; 15'h14B6: d <= 8'hC0; 15'h14B7: d <= 8'hC0;
                15'h14B8: d <= 8'hC0; 15'h14B9: d <= 8'hC0; 15'h14BA: d <= 8'hC0; 15'h14BB: d <= 8'hC0;
                15'h14BC: d <= 8'hC0; 15'h14BD: d <= 8'hC0; 15'h14BE: d <= 8'hC0; 15'h14BF: d <= 8'hC0;
                15'h14C0: d <= 8'hC0; 15'h14C1: d <= 8'hC0; 15'h14C2: d <= 8'hC0; 15'h14C3: d <= 8'hC0;
                15'h14C4: d <= 8'hC0; 15'h14C5: d <= 8'hC0; 15'h14C6: d <= 8'hC0; 15'h14C7: d <= 8'hC0;
                15'h14C8: d <= 8'hC0; 15'h14C9: d <= 8'hC0; 15'h14CA: d <= 8'hC0; 15'h14CB: d <= 8'hC0;
                15'h14CC: d <= 8'hC0; 15'h14CD: d <= 8'hC0; 15'h14CE: d <= 8'hC0; 15'h14CF: d <= 8'hC0;
                15'h14D0: d <= 8'hC0; 15'h14D1: d <= 8'hC0; 15'h14D2: d <= 8'hC0; 15'h14D3: d <= 8'hC0;
                15'h14D4: d <= 8'hC0; 15'h14D5: d <= 8'hC0; 15'h14D6: d <= 8'hC0; 15'h14D7: d <= 8'hC0;
                15'h14D8: d <= 8'hC0; 15'h14D9: d <= 8'hC0; 15'h14DA: d <= 8'hC0; 15'h14DB: d <= 8'hC0;
                15'h14DC: d <= 8'hC0; 15'h14DD: d <= 8'hC0; 15'h14DE: d <= 8'hC0; 15'h14DF: d <= 8'hC0;
                15'h14E0: d <= 8'hC0; 15'h14E1: d <= 8'hC0; 15'h14E2: d <= 8'hC0; 15'h14E3: d <= 8'hC0;
                15'h14E4: d <= 8'hC0; 15'h14E5: d <= 8'hC0; 15'h14E6: d <= 8'hC0; 15'h14E7: d <= 8'hC0;
                15'h14E8: d <= 8'hC0; 15'h14E9: d <= 8'hC0; 15'h14EA: d <= 8'hC0; 15'h14EB: d <= 8'hC0;
                15'h14EC: d <= 8'hC0; 15'h14ED: d <= 8'hC0; 15'h14EE: d <= 8'hC0; 15'h14EF: d <= 8'hC0;
                15'h14F0: d <= 8'hC0; 15'h14F1: d <= 8'hC0; 15'h14F2: d <= 8'hC0; 15'h14F3: d <= 8'hC0;
                15'h14F4: d <= 8'hC0; 15'h14F5: d <= 8'hC0; 15'h14F6: d <= 8'hC0; 15'h14F7: d <= 8'hC0;
                15'h14F8: d <= 8'hC0; 15'h14F9: d <= 8'hC0; 15'h14FA: d <= 8'hC0; 15'h14FB: d <= 8'hC0;
                15'h14FC: d <= 8'hC0; 15'h14FD: d <= 8'hC0; 15'h14FE: d <= 8'hC0; 15'h14FF: d <= 8'hC0;
                15'h1500: d <= 8'hC0; 15'h1501: d <= 8'hC0; 15'h1502: d <= 8'hC0; 15'h1503: d <= 8'hC0;
                15'h1504: d <= 8'hC0; 15'h1505: d <= 8'hC0; 15'h1506: d <= 8'hC0; 15'h1507: d <= 8'hC0;
                15'h1508: d <= 8'hC0; 15'h1509: d <= 8'hC0; 15'h150A: d <= 8'hC0; 15'h150B: d <= 8'hC0;
                15'h150C: d <= 8'hC0; 15'h150D: d <= 8'hC0; 15'h150E: d <= 8'hC0; 15'h150F: d <= 8'hC0;
                15'h1510: d <= 8'hC0; 15'h1511: d <= 8'hC0; 15'h1512: d <= 8'hC0; 15'h1513: d <= 8'hC0;
                15'h1514: d <= 8'hC0; 15'h1515: d <= 8'hC0; 15'h1516: d <= 8'hC0; 15'h1517: d <= 8'hC0;
                15'h1518: d <= 8'hC0; 15'h1519: d <= 8'hC0; 15'h151A: d <= 8'hC0; 15'h151B: d <= 8'hC0;
                15'h151C: d <= 8'hC0; 15'h151D: d <= 8'hC0; 15'h151E: d <= 8'hC0; 15'h151F: d <= 8'hC0;
                15'h1520: d <= 8'hC0; 15'h1521: d <= 8'hC0; 15'h1522: d <= 8'hC0; 15'h1523: d <= 8'hC0;
                15'h1524: d <= 8'hC0; 15'h1525: d <= 8'hC0; 15'h1526: d <= 8'hC0; 15'h1527: d <= 8'hC0;
                15'h1528: d <= 8'hC0; 15'h1529: d <= 8'hC0; 15'h152A: d <= 8'hC0; 15'h152B: d <= 8'hC0;
                15'h152C: d <= 8'hC0; 15'h152D: d <= 8'hC0; 15'h152E: d <= 8'hC0; 15'h152F: d <= 8'hC0;
                15'h1530: d <= 8'hC0; 15'h1531: d <= 8'hC0; 15'h1532: d <= 8'hC0; 15'h1533: d <= 8'hC0;
                15'h1534: d <= 8'hC0; 15'h1535: d <= 8'hC0; 15'h1536: d <= 8'hC0; 15'h1537: d <= 8'hC0;
                15'h1538: d <= 8'hC0; 15'h1539: d <= 8'hC0; 15'h153A: d <= 8'hC0; 15'h153B: d <= 8'hC0;
                15'h153C: d <= 8'hC0; 15'h153D: d <= 8'hC0; 15'h153E: d <= 8'hC0; 15'h153F: d <= 8'hC0;
                15'h1540: d <= 8'hC0; 15'h1541: d <= 8'hC0; 15'h1542: d <= 8'hC0; 15'h1543: d <= 8'hC0;
                15'h1544: d <= 8'hC0; 15'h1545: d <= 8'hC0; 15'h1546: d <= 8'hC0; 15'h1547: d <= 8'hC0;
                15'h1548: d <= 8'hC0; 15'h1549: d <= 8'hC0; 15'h154A: d <= 8'hC0; 15'h154B: d <= 8'hC0;
                15'h154C: d <= 8'hC0; 15'h154D: d <= 8'hC0; 15'h154E: d <= 8'hC0; 15'h154F: d <= 8'hC0;
                15'h1550: d <= 8'hC0; 15'h1551: d <= 8'hC0; 15'h1552: d <= 8'hC0; 15'h1553: d <= 8'hC0;
                15'h1554: d <= 8'hC0; 15'h1555: d <= 8'hC0; 15'h1556: d <= 8'hC0; 15'h1557: d <= 8'hC0;
                15'h1558: d <= 8'hC0; 15'h1559: d <= 8'hC0; 15'h155A: d <= 8'hC0; 15'h155B: d <= 8'hC0;
                15'h155C: d <= 8'hC0; 15'h155D: d <= 8'hC0; 15'h155E: d <= 8'hC0; 15'h155F: d <= 8'hC0;
                15'h1560: d <= 8'hC0; 15'h1561: d <= 8'hC0; 15'h1562: d <= 8'hC0; 15'h1563: d <= 8'hC0;
                15'h1564: d <= 8'hC0; 15'h1565: d <= 8'hC0; 15'h1566: d <= 8'hC0; 15'h1567: d <= 8'hC0;
                15'h1568: d <= 8'hC0; 15'h1569: d <= 8'hC0; 15'h156A: d <= 8'hC0; 15'h156B: d <= 8'hC0;
                15'h156C: d <= 8'hC0; 15'h156D: d <= 8'hC0; 15'h156E: d <= 8'hC0; 15'h156F: d <= 8'hC0;
                15'h1570: d <= 8'hC0; 15'h1571: d <= 8'hC0; 15'h1572: d <= 8'hC0; 15'h1573: d <= 8'hC0;
                15'h1574: d <= 8'hC0; 15'h1575: d <= 8'hC0; 15'h1576: d <= 8'hC0; 15'h1577: d <= 8'hC0;
                15'h1578: d <= 8'hC0; 15'h1579: d <= 8'hC0; 15'h157A: d <= 8'hC0; 15'h157B: d <= 8'hC0;
                15'h157C: d <= 8'hC0; 15'h157D: d <= 8'hC0; 15'h157E: d <= 8'hC0; 15'h157F: d <= 8'hC0;
                15'h1580: d <= 8'hC0; 15'h1581: d <= 8'hC0; 15'h1582: d <= 8'hC0; 15'h1583: d <= 8'hC0;
                15'h1584: d <= 8'hC0; 15'h1585: d <= 8'hC0; 15'h1586: d <= 8'hC0; 15'h1587: d <= 8'hC0;
                15'h1588: d <= 8'hC0; 15'h1589: d <= 8'hC0; 15'h158A: d <= 8'hC0; 15'h158B: d <= 8'hC0;
                15'h158C: d <= 8'hC0; 15'h158D: d <= 8'hC0; 15'h158E: d <= 8'hC0; 15'h158F: d <= 8'hC0;
                15'h1590: d <= 8'hC0; 15'h1591: d <= 8'hC0; 15'h1592: d <= 8'hC0; 15'h1593: d <= 8'hC0;
                15'h1594: d <= 8'hC0; 15'h1595: d <= 8'hC0; 15'h1596: d <= 8'hC0; 15'h1597: d <= 8'hC0;
                15'h1598: d <= 8'hC0; 15'h1599: d <= 8'hC0; 15'h159A: d <= 8'hC0; 15'h159B: d <= 8'hC0;
                15'h159C: d <= 8'hC0; 15'h159D: d <= 8'hC0; 15'h159E: d <= 8'hC0; 15'h159F: d <= 8'hC0;
                15'h15A0: d <= 8'hC0; 15'h15A1: d <= 8'hC0; 15'h15A2: d <= 8'hC0; 15'h15A3: d <= 8'hC0;
                15'h15A4: d <= 8'hC0; 15'h15A5: d <= 8'hC0; 15'h15A6: d <= 8'hC0; 15'h15A7: d <= 8'hC0;
                15'h15A8: d <= 8'hC0; 15'h15A9: d <= 8'hC0; 15'h15AA: d <= 8'hC0; 15'h15AB: d <= 8'hC0;
                15'h15AC: d <= 8'hC0; 15'h15AD: d <= 8'hC0; 15'h15AE: d <= 8'hC0; 15'h15AF: d <= 8'hC0;
                15'h15B0: d <= 8'hC0; 15'h15B1: d <= 8'hC0; 15'h15B2: d <= 8'hC0; 15'h15B3: d <= 8'hC0;
                15'h15B4: d <= 8'hC0; 15'h15B5: d <= 8'hC0; 15'h15B6: d <= 8'hC0; 15'h15B7: d <= 8'hC0;
                15'h15B8: d <= 8'hC0; 15'h15B9: d <= 8'hC0; 15'h15BA: d <= 8'hC0; 15'h15BB: d <= 8'hC0;
                15'h15BC: d <= 8'hC0; 15'h15BD: d <= 8'hC0; 15'h15BE: d <= 8'hC0; 15'h15BF: d <= 8'hC0;
                15'h15C0: d <= 8'hC0; 15'h15C1: d <= 8'hC0; 15'h15C2: d <= 8'hC0; 15'h15C3: d <= 8'hC0;
                15'h15C4: d <= 8'hC0; 15'h15C5: d <= 8'hC0; 15'h15C6: d <= 8'hC0; 15'h15C7: d <= 8'hC0;
                15'h15C8: d <= 8'hC0; 15'h15C9: d <= 8'hC0; 15'h15CA: d <= 8'hC0; 15'h15CB: d <= 8'hC0;
                15'h15CC: d <= 8'hC0; 15'h15CD: d <= 8'hC0; 15'h15CE: d <= 8'hC0; 15'h15CF: d <= 8'hC0;
                15'h15D0: d <= 8'hC0; 15'h15D1: d <= 8'hC0; 15'h15D2: d <= 8'hC0; 15'h15D3: d <= 8'hC0;
                15'h15D4: d <= 8'hC0; 15'h15D5: d <= 8'hC0; 15'h15D6: d <= 8'hC0; 15'h15D7: d <= 8'hC0;
                15'h15D8: d <= 8'hC0; 15'h15D9: d <= 8'hC0; 15'h15DA: d <= 8'hC0; 15'h15DB: d <= 8'hC0;
                15'h15DC: d <= 8'hC0; 15'h15DD: d <= 8'hC0; 15'h15DE: d <= 8'hC0; 15'h15DF: d <= 8'hC0;
                15'h15E0: d <= 8'hC0; 15'h15E1: d <= 8'hC0; 15'h15E2: d <= 8'hC0; 15'h15E3: d <= 8'hC0;
                15'h15E4: d <= 8'hC0; 15'h15E5: d <= 8'hC0; 15'h15E6: d <= 8'hC0; 15'h15E7: d <= 8'hC0;
                15'h15E8: d <= 8'hC0; 15'h15E9: d <= 8'hC0; 15'h15EA: d <= 8'hC0; 15'h15EB: d <= 8'hC0;
                15'h15EC: d <= 8'hC0; 15'h15ED: d <= 8'hC0; 15'h15EE: d <= 8'hC0; 15'h15EF: d <= 8'hC0;
                15'h15F0: d <= 8'hC0; 15'h15F1: d <= 8'hC0; 15'h15F2: d <= 8'hC0; 15'h15F3: d <= 8'hC0;
                15'h15F4: d <= 8'hC0; 15'h15F5: d <= 8'hC0; 15'h15F6: d <= 8'hC0; 15'h15F7: d <= 8'hC0;
                15'h15F8: d <= 8'hC0; 15'h15F9: d <= 8'hC0; 15'h15FA: d <= 8'hC0; 15'h15FB: d <= 8'hC0;
                15'h15FC: d <= 8'hC0; 15'h15FD: d <= 8'hC0; 15'h15FE: d <= 8'hC0; 15'h15FF: d <= 8'hC0;
                15'h1600: d <= 8'hC0; 15'h1601: d <= 8'hC0; 15'h1602: d <= 8'hC0; 15'h1603: d <= 8'hC0;
                15'h1604: d <= 8'hC0; 15'h1605: d <= 8'hC0; 15'h1606: d <= 8'hC0; 15'h1607: d <= 8'hC0;
                15'h1608: d <= 8'hC0; 15'h1609: d <= 8'hC0; 15'h160A: d <= 8'hC0; 15'h160B: d <= 8'hC0;
                15'h160C: d <= 8'hC0; 15'h160D: d <= 8'hC0; 15'h160E: d <= 8'hC0; 15'h160F: d <= 8'hC0;
                15'h1610: d <= 8'hC0; 15'h1611: d <= 8'hC0; 15'h1612: d <= 8'hC0; 15'h1613: d <= 8'hC0;
                15'h1614: d <= 8'hC0; 15'h1615: d <= 8'hC0; 15'h1616: d <= 8'hC0; 15'h1617: d <= 8'hC0;
                15'h1618: d <= 8'hC0; 15'h1619: d <= 8'hC0; 15'h161A: d <= 8'hC0; 15'h161B: d <= 8'hC0;
                15'h161C: d <= 8'hC0; 15'h161D: d <= 8'hC0; 15'h161E: d <= 8'hC0; 15'h161F: d <= 8'hC0;
                15'h1620: d <= 8'hC0; 15'h1621: d <= 8'hC0; 15'h1622: d <= 8'hC0; 15'h1623: d <= 8'hC0;
                15'h1624: d <= 8'hC0; 15'h1625: d <= 8'hC0; 15'h1626: d <= 8'hC0; 15'h1627: d <= 8'hC0;
                15'h1628: d <= 8'hC0; 15'h1629: d <= 8'hC0; 15'h162A: d <= 8'hC0; 15'h162B: d <= 8'hC0;
                15'h162C: d <= 8'hC0; 15'h162D: d <= 8'hC0; 15'h162E: d <= 8'hC0; 15'h162F: d <= 8'hC0;
                15'h1630: d <= 8'hC0; 15'h1631: d <= 8'hC0; 15'h1632: d <= 8'hC0; 15'h1633: d <= 8'hC0;
                15'h1634: d <= 8'hC0; 15'h1635: d <= 8'hC0; 15'h1636: d <= 8'hC0; 15'h1637: d <= 8'hC0;
                15'h1638: d <= 8'hC0; 15'h1639: d <= 8'hC0; 15'h163A: d <= 8'hC0; 15'h163B: d <= 8'hC0;
                15'h163C: d <= 8'hC0; 15'h163D: d <= 8'hC0; 15'h163E: d <= 8'hC0; 15'h163F: d <= 8'hC0;
                15'h1640: d <= 8'hC0; 15'h1641: d <= 8'hC0; 15'h1642: d <= 8'hC0; 15'h1643: d <= 8'hC0;
                15'h1644: d <= 8'hC0; 15'h1645: d <= 8'hC0; 15'h1646: d <= 8'hC0; 15'h1647: d <= 8'hC0;
                15'h1648: d <= 8'hC0; 15'h1649: d <= 8'hC0; 15'h164A: d <= 8'hC0; 15'h164B: d <= 8'hC0;
                15'h164C: d <= 8'hC0; 15'h164D: d <= 8'hC0; 15'h164E: d <= 8'hC0; 15'h164F: d <= 8'hC0;
                15'h1650: d <= 8'hC0; 15'h1651: d <= 8'hC0; 15'h1652: d <= 8'hC0; 15'h1653: d <= 8'hC0;
                15'h1654: d <= 8'hC0; 15'h1655: d <= 8'hC0; 15'h1656: d <= 8'hC0; 15'h1657: d <= 8'hC0;
                15'h1658: d <= 8'hC0; 15'h1659: d <= 8'hC0; 15'h165A: d <= 8'hC0; 15'h165B: d <= 8'hC0;
                15'h165C: d <= 8'hC0; 15'h165D: d <= 8'hC0; 15'h165E: d <= 8'hC0; 15'h165F: d <= 8'hC0;
                15'h1660: d <= 8'hC0; 15'h1661: d <= 8'hC0; 15'h1662: d <= 8'hC0; 15'h1663: d <= 8'hC0;
                15'h1664: d <= 8'hC0; 15'h1665: d <= 8'hC0; 15'h1666: d <= 8'hC0; 15'h1667: d <= 8'hC0;
                15'h1668: d <= 8'hC0; 15'h1669: d <= 8'hC0; 15'h166A: d <= 8'hC0; 15'h166B: d <= 8'hC0;
                15'h166C: d <= 8'hC0; 15'h166D: d <= 8'hC0; 15'h166E: d <= 8'hC0; 15'h166F: d <= 8'hC0;
                15'h1670: d <= 8'hC0; 15'h1671: d <= 8'hC0; 15'h1672: d <= 8'hC0; 15'h1673: d <= 8'hC0;
                15'h1674: d <= 8'hC0; 15'h1675: d <= 8'hC0; 15'h1676: d <= 8'hC0; 15'h1677: d <= 8'hC0;
                15'h1678: d <= 8'hC0; 15'h1679: d <= 8'hC0; 15'h167A: d <= 8'hC0; 15'h167B: d <= 8'hC0;
                15'h167C: d <= 8'hC0; 15'h167D: d <= 8'hC0; 15'h167E: d <= 8'hC0; 15'h167F: d <= 8'hC0;
                15'h1680: d <= 8'hC0; 15'h1681: d <= 8'hC0; 15'h1682: d <= 8'hC0; 15'h1683: d <= 8'hC0;
                15'h1684: d <= 8'hC0; 15'h1685: d <= 8'hC0; 15'h1686: d <= 8'hC0; 15'h1687: d <= 8'hC0;
                15'h1688: d <= 8'hC0; 15'h1689: d <= 8'hC0; 15'h168A: d <= 8'hC0; 15'h168B: d <= 8'hC0;
                15'h168C: d <= 8'hC0; 15'h168D: d <= 8'hC0; 15'h168E: d <= 8'hC0; 15'h168F: d <= 8'hC0;
                15'h1690: d <= 8'hC0; 15'h1691: d <= 8'hC0; 15'h1692: d <= 8'hC0; 15'h1693: d <= 8'hC0;
                15'h1694: d <= 8'hC0; 15'h1695: d <= 8'hC0; 15'h1696: d <= 8'hC0; 15'h1697: d <= 8'hC0;
                15'h1698: d <= 8'hC0; 15'h1699: d <= 8'hC0; 15'h169A: d <= 8'hC0; 15'h169B: d <= 8'hC0;
                15'h169C: d <= 8'hC0; 15'h169D: d <= 8'hC0; 15'h169E: d <= 8'hC0; 15'h169F: d <= 8'hC0;
                15'h16A0: d <= 8'hC0; 15'h16A1: d <= 8'hC0; 15'h16A2: d <= 8'hC0; 15'h16A3: d <= 8'hC0;
                15'h16A4: d <= 8'hC0; 15'h16A5: d <= 8'hC0; 15'h16A6: d <= 8'hC0; 15'h16A7: d <= 8'hC0;
                15'h16A8: d <= 8'hC0; 15'h16A9: d <= 8'hC0; 15'h16AA: d <= 8'hC0; 15'h16AB: d <= 8'hC0;
                15'h16AC: d <= 8'hC0; 15'h16AD: d <= 8'hC0; 15'h16AE: d <= 8'hC0; 15'h16AF: d <= 8'hC0;
                15'h16B0: d <= 8'hC0; 15'h16B1: d <= 8'hC0; 15'h16B2: d <= 8'hC0; 15'h16B3: d <= 8'hC0;
                15'h16B4: d <= 8'hC0; 15'h16B5: d <= 8'hC0; 15'h16B6: d <= 8'hC0; 15'h16B7: d <= 8'hC0;
                15'h16B8: d <= 8'hC0; 15'h16B9: d <= 8'hC0; 15'h16BA: d <= 8'hC0; 15'h16BB: d <= 8'hC0;
                15'h16BC: d <= 8'hC0; 15'h16BD: d <= 8'hC0; 15'h16BE: d <= 8'hC0; 15'h16BF: d <= 8'hC0;
                15'h16C0: d <= 8'hC0; 15'h16C1: d <= 8'hC0; 15'h16C2: d <= 8'hC0; 15'h16C3: d <= 8'hC0;
                15'h16C4: d <= 8'hC0; 15'h16C5: d <= 8'hC0; 15'h16C6: d <= 8'hC0; 15'h16C7: d <= 8'hC0;
                15'h16C8: d <= 8'hC0; 15'h16C9: d <= 8'hC0; 15'h16CA: d <= 8'hC0; 15'h16CB: d <= 8'hC0;
                15'h16CC: d <= 8'hC0; 15'h16CD: d <= 8'hC0; 15'h16CE: d <= 8'hC0; 15'h16CF: d <= 8'hC0;
                15'h16D0: d <= 8'hC0; 15'h16D1: d <= 8'hC0; 15'h16D2: d <= 8'hC0; 15'h16D3: d <= 8'hC0;
                15'h16D4: d <= 8'hC0; 15'h16D5: d <= 8'hC0; 15'h16D6: d <= 8'hC0; 15'h16D7: d <= 8'hC0;
                15'h16D8: d <= 8'hC0; 15'h16D9: d <= 8'hC0; 15'h16DA: d <= 8'hC0; 15'h16DB: d <= 8'hC0;
                15'h16DC: d <= 8'hC0; 15'h16DD: d <= 8'hC0; 15'h16DE: d <= 8'hC0; 15'h16DF: d <= 8'hC0;
                15'h16E0: d <= 8'hC0; 15'h16E1: d <= 8'hC0; 15'h16E2: d <= 8'hC0; 15'h16E3: d <= 8'hC0;
                15'h16E4: d <= 8'hC0; 15'h16E5: d <= 8'hC0; 15'h16E6: d <= 8'hC0; 15'h16E7: d <= 8'hC0;
                15'h16E8: d <= 8'hC0; 15'h16E9: d <= 8'hC0; 15'h16EA: d <= 8'hC0; 15'h16EB: d <= 8'hC0;
                15'h16EC: d <= 8'hC0; 15'h16ED: d <= 8'hC0; 15'h16EE: d <= 8'hC0; 15'h16EF: d <= 8'hC0;
                15'h16F0: d <= 8'hC0; 15'h16F1: d <= 8'hC0; 15'h16F2: d <= 8'hC0; 15'h16F3: d <= 8'hC0;
                15'h16F4: d <= 8'hC0; 15'h16F5: d <= 8'hC0; 15'h16F6: d <= 8'hC0; 15'h16F7: d <= 8'hC0;
                15'h16F8: d <= 8'hC0; 15'h16F9: d <= 8'hC0; 15'h16FA: d <= 8'hC0; 15'h16FB: d <= 8'hC0;
                15'h16FC: d <= 8'hC0; 15'h16FD: d <= 8'hC0; 15'h16FE: d <= 8'hC0; 15'h16FF: d <= 8'hC0;
                15'h1700: d <= 8'hC0; 15'h1701: d <= 8'hC0; 15'h1702: d <= 8'hC0; 15'h1703: d <= 8'hC0;
                15'h1704: d <= 8'hC0; 15'h1705: d <= 8'hC0; 15'h1706: d <= 8'hC0; 15'h1707: d <= 8'hC0;
                15'h1708: d <= 8'hC0; 15'h1709: d <= 8'hC0; 15'h170A: d <= 8'hC0; 15'h170B: d <= 8'hC0;
                15'h170C: d <= 8'hC0; 15'h170D: d <= 8'hC0; 15'h170E: d <= 8'hC0; 15'h170F: d <= 8'hC0;
                15'h1710: d <= 8'hC0; 15'h1711: d <= 8'hC0; 15'h1712: d <= 8'hC0; 15'h1713: d <= 8'hC0;
                15'h1714: d <= 8'hC0; 15'h1715: d <= 8'hC0; 15'h1716: d <= 8'hC0; 15'h1717: d <= 8'hC0;
                15'h1718: d <= 8'hC0; 15'h1719: d <= 8'hC0; 15'h171A: d <= 8'hC0; 15'h171B: d <= 8'hC0;
                15'h171C: d <= 8'hC0; 15'h171D: d <= 8'hC0; 15'h171E: d <= 8'hC0; 15'h171F: d <= 8'hC0;
                15'h1720: d <= 8'hC0; 15'h1721: d <= 8'hC0; 15'h1722: d <= 8'hC0; 15'h1723: d <= 8'hC0;
                15'h1724: d <= 8'hC0; 15'h1725: d <= 8'hC0; 15'h1726: d <= 8'hC0; 15'h1727: d <= 8'hC0;
                15'h1728: d <= 8'hC0; 15'h1729: d <= 8'hC0; 15'h172A: d <= 8'hC0; 15'h172B: d <= 8'hC0;
                15'h172C: d <= 8'hC0; 15'h172D: d <= 8'hC0; 15'h172E: d <= 8'hC0; 15'h172F: d <= 8'hC0;
                15'h1730: d <= 8'hC0; 15'h1731: d <= 8'hC0; 15'h1732: d <= 8'hC0; 15'h1733: d <= 8'hC0;
                15'h1734: d <= 8'hC0; 15'h1735: d <= 8'hC0; 15'h1736: d <= 8'hC0; 15'h1737: d <= 8'hC0;
                15'h1738: d <= 8'hC0; 15'h1739: d <= 8'hC0; 15'h173A: d <= 8'hC0; 15'h173B: d <= 8'hC0;
                15'h173C: d <= 8'hC0; 15'h173D: d <= 8'hC0; 15'h173E: d <= 8'hC0; 15'h173F: d <= 8'hC0;
                15'h1740: d <= 8'hC0; 15'h1741: d <= 8'hC0; 15'h1742: d <= 8'hC0; 15'h1743: d <= 8'hC0;
                15'h1744: d <= 8'hC0; 15'h1745: d <= 8'hC0; 15'h1746: d <= 8'hC0; 15'h1747: d <= 8'hC0;
                15'h1748: d <= 8'hC0; 15'h1749: d <= 8'hC0; 15'h174A: d <= 8'hC0; 15'h174B: d <= 8'hC0;
                15'h174C: d <= 8'hC0; 15'h174D: d <= 8'hC0; 15'h174E: d <= 8'hC0; 15'h174F: d <= 8'hC0;
                15'h1750: d <= 8'hC0; 15'h1751: d <= 8'hC0; 15'h1752: d <= 8'hC0; 15'h1753: d <= 8'hC0;
                15'h1754: d <= 8'hC0; 15'h1755: d <= 8'hC0; 15'h1756: d <= 8'hC0; 15'h1757: d <= 8'hC0;
                15'h1758: d <= 8'hC0; 15'h1759: d <= 8'hC0; 15'h175A: d <= 8'hC0; 15'h175B: d <= 8'hC0;
                15'h175C: d <= 8'hC0; 15'h175D: d <= 8'hC0; 15'h175E: d <= 8'hC0; 15'h175F: d <= 8'hC0;
                15'h1760: d <= 8'hC0; 15'h1761: d <= 8'hC0; 15'h1762: d <= 8'hC0; 15'h1763: d <= 8'hC0;
                15'h1764: d <= 8'hC0; 15'h1765: d <= 8'hC0; 15'h1766: d <= 8'hC0; 15'h1767: d <= 8'hC0;
                15'h1768: d <= 8'hC0; 15'h1769: d <= 8'hC0; 15'h176A: d <= 8'hC0; 15'h176B: d <= 8'hC0;
                15'h176C: d <= 8'hC0; 15'h176D: d <= 8'hC0; 15'h176E: d <= 8'hC0; 15'h176F: d <= 8'hC0;
                15'h1770: d <= 8'hC0; 15'h1771: d <= 8'hC0; 15'h1772: d <= 8'hC0; 15'h1773: d <= 8'hC0;
                15'h1774: d <= 8'hC0; 15'h1775: d <= 8'hC0; 15'h1776: d <= 8'hC0; 15'h1777: d <= 8'hC0;
                15'h1778: d <= 8'hC0; 15'h1779: d <= 8'hC0; 15'h177A: d <= 8'hC0; 15'h177B: d <= 8'hC0;
                15'h177C: d <= 8'hC0; 15'h177D: d <= 8'hC0; 15'h177E: d <= 8'hC0; 15'h177F: d <= 8'hC0;
                15'h1780: d <= 8'hC0; 15'h1781: d <= 8'hC0; 15'h1782: d <= 8'hC0; 15'h1783: d <= 8'hC0;
                15'h1784: d <= 8'hC0; 15'h1785: d <= 8'hC0; 15'h1786: d <= 8'hC0; 15'h1787: d <= 8'hC0;
                15'h1788: d <= 8'hC0; 15'h1789: d <= 8'hC0; 15'h178A: d <= 8'hC0; 15'h178B: d <= 8'hC0;
                15'h178C: d <= 8'hC0; 15'h178D: d <= 8'hC0; 15'h178E: d <= 8'hC0; 15'h178F: d <= 8'hC0;
                15'h1790: d <= 8'hC0; 15'h1791: d <= 8'hC0; 15'h1792: d <= 8'hC0; 15'h1793: d <= 8'hC0;
                15'h1794: d <= 8'hC0; 15'h1795: d <= 8'hC0; 15'h1796: d <= 8'hC0; 15'h1797: d <= 8'hC0;
                15'h1798: d <= 8'hC0; 15'h1799: d <= 8'hC0; 15'h179A: d <= 8'hC0; 15'h179B: d <= 8'hC0;
                15'h179C: d <= 8'hC0; 15'h179D: d <= 8'hC0; 15'h179E: d <= 8'hC0; 15'h179F: d <= 8'hC0;
                15'h17A0: d <= 8'hC0; 15'h17A1: d <= 8'hC0; 15'h17A2: d <= 8'hC0; 15'h17A3: d <= 8'hC0;
                15'h17A4: d <= 8'hC0; 15'h17A5: d <= 8'hC0; 15'h17A6: d <= 8'hC0; 15'h17A7: d <= 8'hC0;
                15'h17A8: d <= 8'hC0; 15'h17A9: d <= 8'hC0; 15'h17AA: d <= 8'hC0; 15'h17AB: d <= 8'hC0;
                15'h17AC: d <= 8'hC0; 15'h17AD: d <= 8'hC0; 15'h17AE: d <= 8'hC0; 15'h17AF: d <= 8'hC0;
                15'h17B0: d <= 8'hC0; 15'h17B1: d <= 8'hC0; 15'h17B2: d <= 8'hC0; 15'h17B3: d <= 8'hC0;
                15'h17B4: d <= 8'hC0; 15'h17B5: d <= 8'hC0; 15'h17B6: d <= 8'hC0; 15'h17B7: d <= 8'hC0;
                15'h17B8: d <= 8'hC0; 15'h17B9: d <= 8'hC0; 15'h17BA: d <= 8'hC0; 15'h17BB: d <= 8'hC0;
                15'h17BC: d <= 8'hC0; 15'h17BD: d <= 8'hC0; 15'h17BE: d <= 8'hC0; 15'h17BF: d <= 8'hC0;
                15'h17C0: d <= 8'hC0; 15'h17C1: d <= 8'hC0; 15'h17C2: d <= 8'hC0; 15'h17C3: d <= 8'hC0;
                15'h17C4: d <= 8'hC0; 15'h17C5: d <= 8'hC0; 15'h17C6: d <= 8'hC0; 15'h17C7: d <= 8'hC0;
                15'h17C8: d <= 8'hC0; 15'h17C9: d <= 8'hC0; 15'h17CA: d <= 8'hC0; 15'h17CB: d <= 8'hC0;
                15'h17CC: d <= 8'hC0; 15'h17CD: d <= 8'hC0; 15'h17CE: d <= 8'hC0; 15'h17CF: d <= 8'hC0;
                15'h17D0: d <= 8'hC0; 15'h17D1: d <= 8'hC0; 15'h17D2: d <= 8'hC0; 15'h17D3: d <= 8'hC0;
                15'h17D4: d <= 8'hC0; 15'h17D5: d <= 8'hC0; 15'h17D6: d <= 8'hC0; 15'h17D7: d <= 8'hC0;
                15'h17D8: d <= 8'hC0; 15'h17D9: d <= 8'hC0; 15'h17DA: d <= 8'hC0; 15'h17DB: d <= 8'hC0;
                15'h17DC: d <= 8'hC0; 15'h17DD: d <= 8'hC0; 15'h17DE: d <= 8'hC0; 15'h17DF: d <= 8'hC0;
                15'h17E0: d <= 8'hC0; 15'h17E1: d <= 8'hC0; 15'h17E2: d <= 8'hC0; 15'h17E3: d <= 8'hC0;
                15'h17E4: d <= 8'hC0; 15'h17E5: d <= 8'hC0; 15'h17E6: d <= 8'hC0; 15'h17E7: d <= 8'hC0;
                15'h17E8: d <= 8'hC0; 15'h17E9: d <= 8'hC0; 15'h17EA: d <= 8'hC0; 15'h17EB: d <= 8'hC0;
                15'h17EC: d <= 8'hC0; 15'h17ED: d <= 8'hC0; 15'h17EE: d <= 8'hC0; 15'h17EF: d <= 8'hC0;
                15'h17F0: d <= 8'hC0; 15'h17F1: d <= 8'hC0; 15'h17F2: d <= 8'hC0; 15'h17F3: d <= 8'hC0;
                15'h17F4: d <= 8'hC0; 15'h17F5: d <= 8'hC0; 15'h17F6: d <= 8'hC0; 15'h17F7: d <= 8'hC0;
                15'h17F8: d <= 8'hC0; 15'h17F9: d <= 8'hC0; 15'h17FA: d <= 8'hC0; 15'h17FB: d <= 8'hC0;
                15'h17FC: d <= 8'hC0; 15'h17FD: d <= 8'hC0; 15'h17FE: d <= 8'hC0; 15'h17FF: d <= 8'hC0;
                15'h1800: d <= 8'hC0; 15'h1801: d <= 8'hC0; 15'h1802: d <= 8'hC0; 15'h1803: d <= 8'hC0;
                15'h1804: d <= 8'hC0; 15'h1805: d <= 8'hC0; 15'h1806: d <= 8'hC0; 15'h1807: d <= 8'hC0;
                15'h1808: d <= 8'hC0; 15'h1809: d <= 8'hC0; 15'h180A: d <= 8'hC0; 15'h180B: d <= 8'hC0;
                15'h180C: d <= 8'hC0; 15'h180D: d <= 8'hC0; 15'h180E: d <= 8'hC0; 15'h180F: d <= 8'hC0;
                15'h1810: d <= 8'hC0; 15'h1811: d <= 8'hC0; 15'h1812: d <= 8'hC0; 15'h1813: d <= 8'hC0;
                15'h1814: d <= 8'hC0; 15'h1815: d <= 8'hC0; 15'h1816: d <= 8'hC0; 15'h1817: d <= 8'hC0;
                15'h1818: d <= 8'hC0; 15'h1819: d <= 8'hC0; 15'h181A: d <= 8'hC0; 15'h181B: d <= 8'hC0;
                15'h181C: d <= 8'hC0; 15'h181D: d <= 8'hC0; 15'h181E: d <= 8'hC0; 15'h181F: d <= 8'hC0;
                15'h1820: d <= 8'hC0; 15'h1821: d <= 8'hC0; 15'h1822: d <= 8'hC0; 15'h1823: d <= 8'hC0;
                15'h1824: d <= 8'hC0; 15'h1825: d <= 8'hC0; 15'h1826: d <= 8'hC0; 15'h1827: d <= 8'hC0;
                15'h1828: d <= 8'hC0; 15'h1829: d <= 8'hC0; 15'h182A: d <= 8'hC0; 15'h182B: d <= 8'hC0;
                15'h182C: d <= 8'hC0; 15'h182D: d <= 8'hC0; 15'h182E: d <= 8'hC0; 15'h182F: d <= 8'hC0;
                15'h1830: d <= 8'hC0; 15'h1831: d <= 8'hC0; 15'h1832: d <= 8'hC0; 15'h1833: d <= 8'hC0;
                15'h1834: d <= 8'hC0; 15'h1835: d <= 8'hC0; 15'h1836: d <= 8'hC0; 15'h1837: d <= 8'hC0;
                15'h1838: d <= 8'hC0; 15'h1839: d <= 8'hC0; 15'h183A: d <= 8'hC0; 15'h183B: d <= 8'hC0;
                15'h183C: d <= 8'hC0; 15'h183D: d <= 8'hC0; 15'h183E: d <= 8'hC0; 15'h183F: d <= 8'hC0;
                15'h1840: d <= 8'hC0; 15'h1841: d <= 8'hC0; 15'h1842: d <= 8'hC0; 15'h1843: d <= 8'hC0;
                15'h1844: d <= 8'hC0; 15'h1845: d <= 8'hC0; 15'h1846: d <= 8'hC0; 15'h1847: d <= 8'hC0;
                15'h1848: d <= 8'hC0; 15'h1849: d <= 8'hC0; 15'h184A: d <= 8'hC0; 15'h184B: d <= 8'hC0;
                15'h184C: d <= 8'hC0; 15'h184D: d <= 8'hC0; 15'h184E: d <= 8'hC0; 15'h184F: d <= 8'hC0;
                15'h1850: d <= 8'hC0; 15'h1851: d <= 8'hC0; 15'h1852: d <= 8'hC0; 15'h1853: d <= 8'hC0;
                15'h1854: d <= 8'hC0; 15'h1855: d <= 8'hC0; 15'h1856: d <= 8'hC0; 15'h1857: d <= 8'hC0;
                15'h1858: d <= 8'hC0; 15'h1859: d <= 8'hC0; 15'h185A: d <= 8'hC0; 15'h185B: d <= 8'hC0;
                15'h185C: d <= 8'hC0; 15'h185D: d <= 8'hC0; 15'h185E: d <= 8'hC0; 15'h185F: d <= 8'hC0;
                15'h1860: d <= 8'hC0; 15'h1861: d <= 8'hC0; 15'h1862: d <= 8'hC0; 15'h1863: d <= 8'hC0;
                15'h1864: d <= 8'hC0; 15'h1865: d <= 8'hC0; 15'h1866: d <= 8'hC0; 15'h1867: d <= 8'hC0;
                15'h1868: d <= 8'hC0; 15'h1869: d <= 8'hC0; 15'h186A: d <= 8'hC0; 15'h186B: d <= 8'hC0;
                15'h186C: d <= 8'hC0; 15'h186D: d <= 8'hC0; 15'h186E: d <= 8'hC0; 15'h186F: d <= 8'hC0;
                15'h1870: d <= 8'hC0; 15'h1871: d <= 8'hC0; 15'h1872: d <= 8'hC0; 15'h1873: d <= 8'hC0;
                15'h1874: d <= 8'hC0; 15'h1875: d <= 8'hC0; 15'h1876: d <= 8'hC0; 15'h1877: d <= 8'hC0;
                15'h1878: d <= 8'hC0; 15'h1879: d <= 8'hC0; 15'h187A: d <= 8'hC0; 15'h187B: d <= 8'hC0;
                15'h187C: d <= 8'hC0; 15'h187D: d <= 8'hC0; 15'h187E: d <= 8'hC0; 15'h187F: d <= 8'hC0;
                15'h1880: d <= 8'hC0; 15'h1881: d <= 8'hC0; 15'h1882: d <= 8'hC0; 15'h1883: d <= 8'hC0;
                15'h1884: d <= 8'hC0; 15'h1885: d <= 8'hC0; 15'h1886: d <= 8'hC0; 15'h1887: d <= 8'hC0;
                15'h1888: d <= 8'hC0; 15'h1889: d <= 8'hC0; 15'h188A: d <= 8'hC0; 15'h188B: d <= 8'hC0;
                15'h188C: d <= 8'hC0; 15'h188D: d <= 8'hC0; 15'h188E: d <= 8'hC0; 15'h188F: d <= 8'hC0;
                15'h1890: d <= 8'hC0; 15'h1891: d <= 8'hC0; 15'h1892: d <= 8'hC0; 15'h1893: d <= 8'hC0;
                15'h1894: d <= 8'hC0; 15'h1895: d <= 8'hC0; 15'h1896: d <= 8'hC0; 15'h1897: d <= 8'hC0;
                15'h1898: d <= 8'hC0; 15'h1899: d <= 8'hC0; 15'h189A: d <= 8'hC0; 15'h189B: d <= 8'hC0;
                15'h189C: d <= 8'hC0; 15'h189D: d <= 8'hC0; 15'h189E: d <= 8'hC0; 15'h189F: d <= 8'hC0;
                15'h18A0: d <= 8'hC0; 15'h18A1: d <= 8'hC0; 15'h18A2: d <= 8'hC0; 15'h18A3: d <= 8'hC0;
                15'h18A4: d <= 8'hC0; 15'h18A5: d <= 8'hC0; 15'h18A6: d <= 8'hC0; 15'h18A7: d <= 8'hC0;
                15'h18A8: d <= 8'hC0; 15'h18A9: d <= 8'hC0; 15'h18AA: d <= 8'hC0; 15'h18AB: d <= 8'hC0;
                15'h18AC: d <= 8'hC0; 15'h18AD: d <= 8'hC0; 15'h18AE: d <= 8'hC0; 15'h18AF: d <= 8'hC0;
                15'h18B0: d <= 8'hC0; 15'h18B1: d <= 8'hC0; 15'h18B2: d <= 8'hC0; 15'h18B3: d <= 8'hC0;
                15'h18B4: d <= 8'hC0; 15'h18B5: d <= 8'hC0; 15'h18B6: d <= 8'hC0; 15'h18B7: d <= 8'hC0;
                15'h18B8: d <= 8'hC0; 15'h18B9: d <= 8'hC0; 15'h18BA: d <= 8'hC0; 15'h18BB: d <= 8'hC0;
                15'h18BC: d <= 8'hC0; 15'h18BD: d <= 8'hC0; 15'h18BE: d <= 8'hC0; 15'h18BF: d <= 8'hC0;
                15'h18C0: d <= 8'hC0; 15'h18C1: d <= 8'hC0; 15'h18C2: d <= 8'hC0; 15'h18C3: d <= 8'hC0;
                15'h18C4: d <= 8'hC0; 15'h18C5: d <= 8'hC0; 15'h18C6: d <= 8'hC0; 15'h18C7: d <= 8'hC0;
                15'h18C8: d <= 8'hC0; 15'h18C9: d <= 8'hC0; 15'h18CA: d <= 8'hC0; 15'h18CB: d <= 8'hC0;
                15'h18CC: d <= 8'hC0; 15'h18CD: d <= 8'hC0; 15'h18CE: d <= 8'hC0; 15'h18CF: d <= 8'hC0;
                15'h18D0: d <= 8'hC0; 15'h18D1: d <= 8'hC0; 15'h18D2: d <= 8'hC0; 15'h18D3: d <= 8'hC0;
                15'h18D4: d <= 8'hC0; 15'h18D5: d <= 8'hC0; 15'h18D6: d <= 8'hC0; 15'h18D7: d <= 8'hC0;
                15'h18D8: d <= 8'hC0; 15'h18D9: d <= 8'hC0; 15'h18DA: d <= 8'hC0; 15'h18DB: d <= 8'hC0;
                15'h18DC: d <= 8'hC0; 15'h18DD: d <= 8'hC0; 15'h18DE: d <= 8'hC0; 15'h18DF: d <= 8'hC0;
                15'h18E0: d <= 8'hC0; 15'h18E1: d <= 8'hC0; 15'h18E2: d <= 8'hC0; 15'h18E3: d <= 8'hC0;
                15'h18E4: d <= 8'hC0; 15'h18E5: d <= 8'hC0; 15'h18E6: d <= 8'hC0; 15'h18E7: d <= 8'hC0;
                15'h18E8: d <= 8'hC0; 15'h18E9: d <= 8'hC0; 15'h18EA: d <= 8'hC0; 15'h18EB: d <= 8'hC0;
                15'h18EC: d <= 8'hC0; 15'h18ED: d <= 8'hC0; 15'h18EE: d <= 8'hC0; 15'h18EF: d <= 8'hC0;
                15'h18F0: d <= 8'hC0; 15'h18F1: d <= 8'hC0; 15'h18F2: d <= 8'hC0; 15'h18F3: d <= 8'hC0;
                15'h18F4: d <= 8'hC0; 15'h18F5: d <= 8'hC0; 15'h18F6: d <= 8'hC0; 15'h18F7: d <= 8'hC0;
                15'h18F8: d <= 8'hC0; 15'h18F9: d <= 8'hC0; 15'h18FA: d <= 8'hC0; 15'h18FB: d <= 8'hC0;
                15'h18FC: d <= 8'hC0; 15'h18FD: d <= 8'hC0; 15'h18FE: d <= 8'hC0; 15'h18FF: d <= 8'hC0;
                15'h1900: d <= 8'hC0; 15'h1901: d <= 8'hC0; 15'h1902: d <= 8'hC0; 15'h1903: d <= 8'hC0;
                15'h1904: d <= 8'hC0; 15'h1905: d <= 8'hC0; 15'h1906: d <= 8'hC0; 15'h1907: d <= 8'hC0;
                15'h1908: d <= 8'hC0; 15'h1909: d <= 8'hC0; 15'h190A: d <= 8'hC0; 15'h190B: d <= 8'hC0;
                15'h190C: d <= 8'hC0; 15'h190D: d <= 8'hC0; 15'h190E: d <= 8'hC0; 15'h190F: d <= 8'hC0;
                15'h1910: d <= 8'hC0; 15'h1911: d <= 8'hC0; 15'h1912: d <= 8'hC0; 15'h1913: d <= 8'hC0;
                15'h1914: d <= 8'hC0; 15'h1915: d <= 8'hC0; 15'h1916: d <= 8'hC0; 15'h1917: d <= 8'hC0;
                15'h1918: d <= 8'hC0; 15'h1919: d <= 8'hC0; 15'h191A: d <= 8'hC0; 15'h191B: d <= 8'hC0;
                15'h191C: d <= 8'hC0; 15'h191D: d <= 8'hC0; 15'h191E: d <= 8'hC0; 15'h191F: d <= 8'hC0;
                15'h1920: d <= 8'hC0; 15'h1921: d <= 8'hC0; 15'h1922: d <= 8'hC0; 15'h1923: d <= 8'hC0;
                15'h1924: d <= 8'hC0; 15'h1925: d <= 8'hC0; 15'h1926: d <= 8'hC0; 15'h1927: d <= 8'hC0;
                15'h1928: d <= 8'hC0; 15'h1929: d <= 8'hC0; 15'h192A: d <= 8'hC0; 15'h192B: d <= 8'hC0;
                15'h192C: d <= 8'hC0; 15'h192D: d <= 8'hC0; 15'h192E: d <= 8'hC0; 15'h192F: d <= 8'hC0;
                15'h1930: d <= 8'hC0; 15'h1931: d <= 8'hC0; 15'h1932: d <= 8'hC0; 15'h1933: d <= 8'hC0;
                15'h1934: d <= 8'hC0; 15'h1935: d <= 8'hC0; 15'h1936: d <= 8'hC0; 15'h1937: d <= 8'hC0;
                15'h1938: d <= 8'hC0; 15'h1939: d <= 8'hC0; 15'h193A: d <= 8'hC0; 15'h193B: d <= 8'hC0;
                15'h193C: d <= 8'hC0; 15'h193D: d <= 8'hC0; 15'h193E: d <= 8'hC0; 15'h193F: d <= 8'hC0;
                15'h1940: d <= 8'hC0; 15'h1941: d <= 8'hC0; 15'h1942: d <= 8'hC0; 15'h1943: d <= 8'hC0;
                15'h1944: d <= 8'hC0; 15'h1945: d <= 8'hC0; 15'h1946: d <= 8'hC0; 15'h1947: d <= 8'hC0;
                15'h1948: d <= 8'hC0; 15'h1949: d <= 8'hC0; 15'h194A: d <= 8'hC0; 15'h194B: d <= 8'hC0;
                15'h194C: d <= 8'hC0; 15'h194D: d <= 8'hC0; 15'h194E: d <= 8'hC0; 15'h194F: d <= 8'hC0;
                15'h1950: d <= 8'hC0; 15'h1951: d <= 8'hC0; 15'h1952: d <= 8'hC0; 15'h1953: d <= 8'hC0;
                15'h1954: d <= 8'hC0; 15'h1955: d <= 8'hC0; 15'h1956: d <= 8'hC0; 15'h1957: d <= 8'hC0;
                15'h1958: d <= 8'hC0; 15'h1959: d <= 8'hC0; 15'h195A: d <= 8'hC0; 15'h195B: d <= 8'hC0;
                15'h195C: d <= 8'hC0; 15'h195D: d <= 8'hC0; 15'h195E: d <= 8'hC0; 15'h195F: d <= 8'hC0;
                15'h1960: d <= 8'hC0; 15'h1961: d <= 8'hC0; 15'h1962: d <= 8'hC0; 15'h1963: d <= 8'hC0;
                15'h1964: d <= 8'hC0; 15'h1965: d <= 8'hC0; 15'h1966: d <= 8'hC0; 15'h1967: d <= 8'hC0;
                15'h1968: d <= 8'hC0; 15'h1969: d <= 8'hC0; 15'h196A: d <= 8'hC0; 15'h196B: d <= 8'hC0;
                15'h196C: d <= 8'hC0; 15'h196D: d <= 8'hC0; 15'h196E: d <= 8'hC0; 15'h196F: d <= 8'hC0;
                15'h1970: d <= 8'hC0; 15'h1971: d <= 8'hC0; 15'h1972: d <= 8'hC0; 15'h1973: d <= 8'hC0;
                15'h1974: d <= 8'hC0; 15'h1975: d <= 8'hC0; 15'h1976: d <= 8'hC0; 15'h1977: d <= 8'hC0;
                15'h1978: d <= 8'hC0; 15'h1979: d <= 8'hC0; 15'h197A: d <= 8'hC0; 15'h197B: d <= 8'hC0;
                15'h197C: d <= 8'hC0; 15'h197D: d <= 8'hC0; 15'h197E: d <= 8'hC0; 15'h197F: d <= 8'hC0;
                15'h1980: d <= 8'hC0; 15'h1981: d <= 8'hC0; 15'h1982: d <= 8'hC0; 15'h1983: d <= 8'hC0;
                15'h1984: d <= 8'hC0; 15'h1985: d <= 8'hC0; 15'h1986: d <= 8'hC0; 15'h1987: d <= 8'hC0;
                15'h1988: d <= 8'hC0; 15'h1989: d <= 8'hC0; 15'h198A: d <= 8'hC0; 15'h198B: d <= 8'hC0;
                15'h198C: d <= 8'hC0; 15'h198D: d <= 8'hC0; 15'h198E: d <= 8'hC0; 15'h198F: d <= 8'hC0;
                15'h1990: d <= 8'hC0; 15'h1991: d <= 8'hC0; 15'h1992: d <= 8'hC0; 15'h1993: d <= 8'hC0;
                15'h1994: d <= 8'hC0; 15'h1995: d <= 8'hC0; 15'h1996: d <= 8'hC0; 15'h1997: d <= 8'hC0;
                15'h1998: d <= 8'hC0; 15'h1999: d <= 8'hC0; 15'h199A: d <= 8'hC0; 15'h199B: d <= 8'hC0;
                15'h199C: d <= 8'hC0; 15'h199D: d <= 8'hC0; 15'h199E: d <= 8'hC0; 15'h199F: d <= 8'hC0;
                15'h19A0: d <= 8'hC0; 15'h19A1: d <= 8'hC0; 15'h19A2: d <= 8'hC0; 15'h19A3: d <= 8'hC0;
                15'h19A4: d <= 8'hC0; 15'h19A5: d <= 8'hC0; 15'h19A6: d <= 8'hC0; 15'h19A7: d <= 8'hC0;
                15'h19A8: d <= 8'hC0; 15'h19A9: d <= 8'hC0; 15'h19AA: d <= 8'hC0; 15'h19AB: d <= 8'hC0;
                15'h19AC: d <= 8'hC0; 15'h19AD: d <= 8'hC0; 15'h19AE: d <= 8'hC0; 15'h19AF: d <= 8'hC0;
                15'h19B0: d <= 8'hC0; 15'h19B1: d <= 8'hC0; 15'h19B2: d <= 8'hC0; 15'h19B3: d <= 8'hC0;
                15'h19B4: d <= 8'hC0; 15'h19B5: d <= 8'hC0; 15'h19B6: d <= 8'hC0; 15'h19B7: d <= 8'hC0;
                15'h19B8: d <= 8'hC0; 15'h19B9: d <= 8'hC0; 15'h19BA: d <= 8'hC0; 15'h19BB: d <= 8'hC0;
                15'h19BC: d <= 8'hC0; 15'h19BD: d <= 8'hC0; 15'h19BE: d <= 8'hC0; 15'h19BF: d <= 8'hC0;
                15'h19C0: d <= 8'hC0; 15'h19C1: d <= 8'hC0; 15'h19C2: d <= 8'hC0; 15'h19C3: d <= 8'hC0;
                15'h19C4: d <= 8'hC0; 15'h19C5: d <= 8'hC0; 15'h19C6: d <= 8'hC0; 15'h19C7: d <= 8'hC0;
                15'h19C8: d <= 8'hC0; 15'h19C9: d <= 8'hC0; 15'h19CA: d <= 8'hC0; 15'h19CB: d <= 8'hC0;
                15'h19CC: d <= 8'hC0; 15'h19CD: d <= 8'hC0; 15'h19CE: d <= 8'hC0; 15'h19CF: d <= 8'hC0;
                15'h19D0: d <= 8'hC0; 15'h19D1: d <= 8'hC0; 15'h19D2: d <= 8'hC0; 15'h19D3: d <= 8'hC0;
                15'h19D4: d <= 8'hC0; 15'h19D5: d <= 8'hC0; 15'h19D6: d <= 8'hC0; 15'h19D7: d <= 8'hC0;
                15'h19D8: d <= 8'hC0; 15'h19D9: d <= 8'hC0; 15'h19DA: d <= 8'hC0; 15'h19DB: d <= 8'hC0;
                15'h19DC: d <= 8'hC0; 15'h19DD: d <= 8'hC0; 15'h19DE: d <= 8'hC0; 15'h19DF: d <= 8'hC0;
                15'h19E0: d <= 8'hC0; 15'h19E1: d <= 8'hC0; 15'h19E2: d <= 8'hC0; 15'h19E3: d <= 8'hC0;
                15'h19E4: d <= 8'hC0; 15'h19E5: d <= 8'hC0; 15'h19E6: d <= 8'hC0; 15'h19E7: d <= 8'hC0;
                15'h19E8: d <= 8'hC0; 15'h19E9: d <= 8'hC0; 15'h19EA: d <= 8'hC0; 15'h19EB: d <= 8'hC0;
                15'h19EC: d <= 8'hC0; 15'h19ED: d <= 8'hC0; 15'h19EE: d <= 8'hC0; 15'h19EF: d <= 8'hC0;
                15'h19F0: d <= 8'hC0; 15'h19F1: d <= 8'hC0; 15'h19F2: d <= 8'hC0; 15'h19F3: d <= 8'hC0;
                15'h19F4: d <= 8'hC0; 15'h19F5: d <= 8'hC0; 15'h19F6: d <= 8'hC0; 15'h19F7: d <= 8'hC0;
                15'h19F8: d <= 8'hC0; 15'h19F9: d <= 8'hC0; 15'h19FA: d <= 8'hC0; 15'h19FB: d <= 8'hC0;
                15'h19FC: d <= 8'hC0; 15'h19FD: d <= 8'hC0; 15'h19FE: d <= 8'hC0; 15'h19FF: d <= 8'hC0;
                15'h1A00: d <= 8'hC0; 15'h1A01: d <= 8'hC0; 15'h1A02: d <= 8'hC0; 15'h1A03: d <= 8'hC0;
                15'h1A04: d <= 8'hC0; 15'h1A05: d <= 8'hC0; 15'h1A06: d <= 8'hC0; 15'h1A07: d <= 8'hC0;
                15'h1A08: d <= 8'hC0; 15'h1A09: d <= 8'hC0; 15'h1A0A: d <= 8'hC0; 15'h1A0B: d <= 8'hC0;
                15'h1A0C: d <= 8'hC0; 15'h1A0D: d <= 8'hC0; 15'h1A0E: d <= 8'hC0; 15'h1A0F: d <= 8'hC0;
                15'h1A10: d <= 8'hC0; 15'h1A11: d <= 8'hC0; 15'h1A12: d <= 8'hC0; 15'h1A13: d <= 8'hC0;
                15'h1A14: d <= 8'hC0; 15'h1A15: d <= 8'hC0; 15'h1A16: d <= 8'hC0; 15'h1A17: d <= 8'hC0;
                15'h1A18: d <= 8'hC0; 15'h1A19: d <= 8'hC0; 15'h1A1A: d <= 8'hC0; 15'h1A1B: d <= 8'hC0;
                15'h1A1C: d <= 8'hC0; 15'h1A1D: d <= 8'hC0; 15'h1A1E: d <= 8'hC0; 15'h1A1F: d <= 8'hC0;
                15'h1A20: d <= 8'hC0; 15'h1A21: d <= 8'hC0; 15'h1A22: d <= 8'hC0; 15'h1A23: d <= 8'hC0;
                15'h1A24: d <= 8'hC0; 15'h1A25: d <= 8'hC0; 15'h1A26: d <= 8'hC0; 15'h1A27: d <= 8'hC0;
                15'h1A28: d <= 8'hC0; 15'h1A29: d <= 8'hC0; 15'h1A2A: d <= 8'hC0; 15'h1A2B: d <= 8'hC0;
                15'h1A2C: d <= 8'hC0; 15'h1A2D: d <= 8'hC0; 15'h1A2E: d <= 8'hC0; 15'h1A2F: d <= 8'hC0;
                15'h1A30: d <= 8'hC0; 15'h1A31: d <= 8'hC0; 15'h1A32: d <= 8'hC0; 15'h1A33: d <= 8'hC0;
                15'h1A34: d <= 8'hC0; 15'h1A35: d <= 8'hC0; 15'h1A36: d <= 8'hC0; 15'h1A37: d <= 8'hC0;
                15'h1A38: d <= 8'hC0; 15'h1A39: d <= 8'hC0; 15'h1A3A: d <= 8'hC0; 15'h1A3B: d <= 8'hC0;
                15'h1A3C: d <= 8'hC0; 15'h1A3D: d <= 8'hC0; 15'h1A3E: d <= 8'hC0; 15'h1A3F: d <= 8'hC0;
                15'h1A40: d <= 8'hC0; 15'h1A41: d <= 8'hC0; 15'h1A42: d <= 8'hC0; 15'h1A43: d <= 8'hC0;
                15'h1A44: d <= 8'hC0; 15'h1A45: d <= 8'hC0; 15'h1A46: d <= 8'hC0; 15'h1A47: d <= 8'hC0;
                15'h1A48: d <= 8'hC0; 15'h1A49: d <= 8'hC0; 15'h1A4A: d <= 8'hC0; 15'h1A4B: d <= 8'hC0;
                15'h1A4C: d <= 8'hC0; 15'h1A4D: d <= 8'hC0; 15'h1A4E: d <= 8'hC0; 15'h1A4F: d <= 8'hC0;
                15'h1A50: d <= 8'hC0; 15'h1A51: d <= 8'hC0; 15'h1A52: d <= 8'hC0; 15'h1A53: d <= 8'hC0;
                15'h1A54: d <= 8'hC0; 15'h1A55: d <= 8'hC0; 15'h1A56: d <= 8'hC0; 15'h1A57: d <= 8'hC0;
                15'h1A58: d <= 8'hC0; 15'h1A59: d <= 8'hC0; 15'h1A5A: d <= 8'hC0; 15'h1A5B: d <= 8'hC0;
                15'h1A5C: d <= 8'hC0; 15'h1A5D: d <= 8'hC0; 15'h1A5E: d <= 8'hC0; 15'h1A5F: d <= 8'hC0;
                15'h1A60: d <= 8'hC0; 15'h1A61: d <= 8'hC0; 15'h1A62: d <= 8'hC0; 15'h1A63: d <= 8'hC0;
                15'h1A64: d <= 8'hC0; 15'h1A65: d <= 8'hC0; 15'h1A66: d <= 8'hC0; 15'h1A67: d <= 8'hC0;
                15'h1A68: d <= 8'hC0; 15'h1A69: d <= 8'hC0; 15'h1A6A: d <= 8'hC0; 15'h1A6B: d <= 8'hC0;
                15'h1A6C: d <= 8'hC0; 15'h1A6D: d <= 8'hC0; 15'h1A6E: d <= 8'hC0; 15'h1A6F: d <= 8'hC0;
                15'h1A70: d <= 8'hC0; 15'h1A71: d <= 8'hC0; 15'h1A72: d <= 8'hC0; 15'h1A73: d <= 8'hC0;
                15'h1A74: d <= 8'hC0; 15'h1A75: d <= 8'hC0; 15'h1A76: d <= 8'hC0; 15'h1A77: d <= 8'hC0;
                15'h1A78: d <= 8'hC0; 15'h1A79: d <= 8'hC0; 15'h1A7A: d <= 8'hC0; 15'h1A7B: d <= 8'hC0;
                15'h1A7C: d <= 8'hC0; 15'h1A7D: d <= 8'hC0; 15'h1A7E: d <= 8'hC0; 15'h1A7F: d <= 8'hC0;
                15'h1A80: d <= 8'hC0; 15'h1A81: d <= 8'hC0; 15'h1A82: d <= 8'hC0; 15'h1A83: d <= 8'hC0;
                15'h1A84: d <= 8'hC0; 15'h1A85: d <= 8'hC0; 15'h1A86: d <= 8'hC0; 15'h1A87: d <= 8'hC0;
                15'h1A88: d <= 8'hC0; 15'h1A89: d <= 8'hC0; 15'h1A8A: d <= 8'hC0; 15'h1A8B: d <= 8'hC0;
                15'h1A8C: d <= 8'hC0; 15'h1A8D: d <= 8'hC0; 15'h1A8E: d <= 8'hC0; 15'h1A8F: d <= 8'hC0;
                15'h1A90: d <= 8'hC0; 15'h1A91: d <= 8'hC0; 15'h1A92: d <= 8'hC0; 15'h1A93: d <= 8'hC0;
                15'h1A94: d <= 8'hC0; 15'h1A95: d <= 8'hC0; 15'h1A96: d <= 8'hC0; 15'h1A97: d <= 8'hC0;
                15'h1A98: d <= 8'hC0; 15'h1A99: d <= 8'hC0; 15'h1A9A: d <= 8'hC0; 15'h1A9B: d <= 8'hC0;
                15'h1A9C: d <= 8'hC0; 15'h1A9D: d <= 8'hC0; 15'h1A9E: d <= 8'hC0; 15'h1A9F: d <= 8'hC0;
                15'h1AA0: d <= 8'hC0; 15'h1AA1: d <= 8'hC0; 15'h1AA2: d <= 8'hC0; 15'h1AA3: d <= 8'hC0;
                15'h1AA4: d <= 8'hC0; 15'h1AA5: d <= 8'hC0; 15'h1AA6: d <= 8'hC0; 15'h1AA7: d <= 8'hC0;
                15'h1AA8: d <= 8'hC0; 15'h1AA9: d <= 8'hC0; 15'h1AAA: d <= 8'hC0; 15'h1AAB: d <= 8'hC0;
                15'h1AAC: d <= 8'hC0; 15'h1AAD: d <= 8'hC0; 15'h1AAE: d <= 8'hC0; 15'h1AAF: d <= 8'hC0;
                15'h1AB0: d <= 8'hC0; 15'h1AB1: d <= 8'hC0; 15'h1AB2: d <= 8'hC0; 15'h1AB3: d <= 8'hC0;
                15'h1AB4: d <= 8'hC0; 15'h1AB5: d <= 8'hC0; 15'h1AB6: d <= 8'hC0; 15'h1AB7: d <= 8'hC0;
                15'h1AB8: d <= 8'hC0; 15'h1AB9: d <= 8'hC0; 15'h1ABA: d <= 8'hC0; 15'h1ABB: d <= 8'hC0;
                15'h1ABC: d <= 8'hC0; 15'h1ABD: d <= 8'hC0; 15'h1ABE: d <= 8'hC0; 15'h1ABF: d <= 8'hC0;
                15'h1AC0: d <= 8'hC0; 15'h1AC1: d <= 8'hC0; 15'h1AC2: d <= 8'hC0; 15'h1AC3: d <= 8'hC0;
                15'h1AC4: d <= 8'hC0; 15'h1AC5: d <= 8'hC0; 15'h1AC6: d <= 8'hC0; 15'h1AC7: d <= 8'hC0;
                15'h1AC8: d <= 8'hC0; 15'h1AC9: d <= 8'hC0; 15'h1ACA: d <= 8'hC0; 15'h1ACB: d <= 8'hC0;
                15'h1ACC: d <= 8'hC0; 15'h1ACD: d <= 8'hC0; 15'h1ACE: d <= 8'hC0; 15'h1ACF: d <= 8'hC0;
                15'h1AD0: d <= 8'hC0; 15'h1AD1: d <= 8'hC0; 15'h1AD2: d <= 8'hC0; 15'h1AD3: d <= 8'hC0;
                15'h1AD4: d <= 8'hC0; 15'h1AD5: d <= 8'hC0; 15'h1AD6: d <= 8'hC0; 15'h1AD7: d <= 8'hC0;
                15'h1AD8: d <= 8'hC0; 15'h1AD9: d <= 8'hC0; 15'h1ADA: d <= 8'hC0; 15'h1ADB: d <= 8'hC0;
                15'h1ADC: d <= 8'hC0; 15'h1ADD: d <= 8'hC0; 15'h1ADE: d <= 8'hC0; 15'h1ADF: d <= 8'hC0;
                15'h1AE0: d <= 8'hC0; 15'h1AE1: d <= 8'hC0; 15'h1AE2: d <= 8'hC0; 15'h1AE3: d <= 8'hC0;
                15'h1AE4: d <= 8'hC0; 15'h1AE5: d <= 8'hC0; 15'h1AE6: d <= 8'hC0; 15'h1AE7: d <= 8'hC0;
                15'h1AE8: d <= 8'hC0; 15'h1AE9: d <= 8'hC0; 15'h1AEA: d <= 8'hC0; 15'h1AEB: d <= 8'hC0;
                15'h1AEC: d <= 8'hC0; 15'h1AED: d <= 8'hC0; 15'h1AEE: d <= 8'hC0; 15'h1AEF: d <= 8'hC0;
                15'h1AF0: d <= 8'hC0; 15'h1AF1: d <= 8'hC0; 15'h1AF2: d <= 8'hC0; 15'h1AF3: d <= 8'hC0;
                15'h1AF4: d <= 8'hC0; 15'h1AF5: d <= 8'hC0; 15'h1AF6: d <= 8'hC0; 15'h1AF7: d <= 8'hC0;
                15'h1AF8: d <= 8'hC0; 15'h1AF9: d <= 8'hC0; 15'h1AFA: d <= 8'hC0; 15'h1AFB: d <= 8'hC0;
                15'h1AFC: d <= 8'hC0; 15'h1AFD: d <= 8'hC0; 15'h1AFE: d <= 8'hC0; 15'h1AFF: d <= 8'hC0;
                15'h1B00: d <= 8'hC0; 15'h1B01: d <= 8'hC0; 15'h1B02: d <= 8'hC0; 15'h1B03: d <= 8'hC0;
                15'h1B04: d <= 8'hC0; 15'h1B05: d <= 8'hC0; 15'h1B06: d <= 8'hC0; 15'h1B07: d <= 8'hC0;
                15'h1B08: d <= 8'hC0; 15'h1B09: d <= 8'hC0; 15'h1B0A: d <= 8'hC0; 15'h1B0B: d <= 8'hC0;
                15'h1B0C: d <= 8'hC0; 15'h1B0D: d <= 8'hC0; 15'h1B0E: d <= 8'hC0; 15'h1B0F: d <= 8'hC0;
                15'h1B10: d <= 8'hC0; 15'h1B11: d <= 8'hC0; 15'h1B12: d <= 8'hC0; 15'h1B13: d <= 8'hC0;
                15'h1B14: d <= 8'hC0; 15'h1B15: d <= 8'hC0; 15'h1B16: d <= 8'hC0; 15'h1B17: d <= 8'hC0;
                15'h1B18: d <= 8'hC0; 15'h1B19: d <= 8'hC0; 15'h1B1A: d <= 8'hC0; 15'h1B1B: d <= 8'hC0;
                15'h1B1C: d <= 8'hC0; 15'h1B1D: d <= 8'hC0; 15'h1B1E: d <= 8'hC0; 15'h1B1F: d <= 8'hC0;
                15'h1B20: d <= 8'hC0; 15'h1B21: d <= 8'hC0; 15'h1B22: d <= 8'hC0; 15'h1B23: d <= 8'hC0;
                15'h1B24: d <= 8'hC0; 15'h1B25: d <= 8'hC0; 15'h1B26: d <= 8'hC0; 15'h1B27: d <= 8'hC0;
                15'h1B28: d <= 8'hC0; 15'h1B29: d <= 8'hC0; 15'h1B2A: d <= 8'hC0; 15'h1B2B: d <= 8'hC0;
                15'h1B2C: d <= 8'hC0; 15'h1B2D: d <= 8'hC0; 15'h1B2E: d <= 8'hC0; 15'h1B2F: d <= 8'hC0;
                15'h1B30: d <= 8'hC0; 15'h1B31: d <= 8'hC0; 15'h1B32: d <= 8'hC0; 15'h1B33: d <= 8'hC0;
                15'h1B34: d <= 8'hC0; 15'h1B35: d <= 8'hC0; 15'h1B36: d <= 8'hC0; 15'h1B37: d <= 8'hC0;
                15'h1B38: d <= 8'hC0; 15'h1B39: d <= 8'hC0; 15'h1B3A: d <= 8'hC0; 15'h1B3B: d <= 8'hC0;
                15'h1B3C: d <= 8'hC0; 15'h1B3D: d <= 8'hC0; 15'h1B3E: d <= 8'hC0; 15'h1B3F: d <= 8'hC0;
                15'h1B40: d <= 8'hC0; 15'h1B41: d <= 8'hC0; 15'h1B42: d <= 8'hC0; 15'h1B43: d <= 8'hC0;
                15'h1B44: d <= 8'hC0; 15'h1B45: d <= 8'hC0; 15'h1B46: d <= 8'hC0; 15'h1B47: d <= 8'hC0;
                15'h1B48: d <= 8'hC0; 15'h1B49: d <= 8'hC0; 15'h1B4A: d <= 8'hC0; 15'h1B4B: d <= 8'hC0;
                15'h1B4C: d <= 8'hC0; 15'h1B4D: d <= 8'hC0; 15'h1B4E: d <= 8'hC0; 15'h1B4F: d <= 8'hC0;
                15'h1B50: d <= 8'hC0; 15'h1B51: d <= 8'hC0; 15'h1B52: d <= 8'hC0; 15'h1B53: d <= 8'hC0;
                15'h1B54: d <= 8'hC0; 15'h1B55: d <= 8'hC0; 15'h1B56: d <= 8'hC0; 15'h1B57: d <= 8'hC0;
                15'h1B58: d <= 8'hC0; 15'h1B59: d <= 8'hC0; 15'h1B5A: d <= 8'hC0; 15'h1B5B: d <= 8'hC0;
                15'h1B5C: d <= 8'hC0; 15'h1B5D: d <= 8'hC0; 15'h1B5E: d <= 8'hC0; 15'h1B5F: d <= 8'hC0;
                15'h1B60: d <= 8'hC0; 15'h1B61: d <= 8'hC0; 15'h1B62: d <= 8'hC0; 15'h1B63: d <= 8'hC0;
                15'h1B64: d <= 8'hC0; 15'h1B65: d <= 8'hC0; 15'h1B66: d <= 8'hC0; 15'h1B67: d <= 8'hC0;
                15'h1B68: d <= 8'hC0; 15'h1B69: d <= 8'hC0; 15'h1B6A: d <= 8'hC0; 15'h1B6B: d <= 8'hC0;
                15'h1B6C: d <= 8'hC0; 15'h1B6D: d <= 8'hC0; 15'h1B6E: d <= 8'hC0; 15'h1B6F: d <= 8'hC0;
                15'h1B70: d <= 8'hC0; 15'h1B71: d <= 8'hC0; 15'h1B72: d <= 8'hC0; 15'h1B73: d <= 8'hC0;
                15'h1B74: d <= 8'hC0; 15'h1B75: d <= 8'hC0; 15'h1B76: d <= 8'hC0; 15'h1B77: d <= 8'hC0;
                15'h1B78: d <= 8'hC0; 15'h1B79: d <= 8'hC0; 15'h1B7A: d <= 8'hC0; 15'h1B7B: d <= 8'hC0;
                15'h1B7C: d <= 8'hC0; 15'h1B7D: d <= 8'hC0; 15'h1B7E: d <= 8'hC0; 15'h1B7F: d <= 8'hC0;
                15'h1B80: d <= 8'hC0; 15'h1B81: d <= 8'hC0; 15'h1B82: d <= 8'hC0; 15'h1B83: d <= 8'hC0;
                15'h1B84: d <= 8'hC0; 15'h1B85: d <= 8'hC0; 15'h1B86: d <= 8'hC0; 15'h1B87: d <= 8'hC0;
                15'h1B88: d <= 8'hC0; 15'h1B89: d <= 8'hC0; 15'h1B8A: d <= 8'hC0; 15'h1B8B: d <= 8'hC0;
                15'h1B8C: d <= 8'hC0; 15'h1B8D: d <= 8'hC0; 15'h1B8E: d <= 8'hC0; 15'h1B8F: d <= 8'hC0;
                15'h1B90: d <= 8'hC0; 15'h1B91: d <= 8'hC0; 15'h1B92: d <= 8'hC0; 15'h1B93: d <= 8'hC0;
                15'h1B94: d <= 8'hC0; 15'h1B95: d <= 8'hC0; 15'h1B96: d <= 8'hC0; 15'h1B97: d <= 8'hC0;
                15'h1B98: d <= 8'hC0; 15'h1B99: d <= 8'hC0; 15'h1B9A: d <= 8'hC0; 15'h1B9B: d <= 8'hC0;
                15'h1B9C: d <= 8'hC0; 15'h1B9D: d <= 8'hC0; 15'h1B9E: d <= 8'hC0; 15'h1B9F: d <= 8'hC0;
                15'h1BA0: d <= 8'hC0; 15'h1BA1: d <= 8'hC0; 15'h1BA2: d <= 8'hC0; 15'h1BA3: d <= 8'hC0;
                15'h1BA4: d <= 8'hC0; 15'h1BA5: d <= 8'hC0; 15'h1BA6: d <= 8'hC0; 15'h1BA7: d <= 8'hC0;
                15'h1BA8: d <= 8'hC0; 15'h1BA9: d <= 8'hC0; 15'h1BAA: d <= 8'hC0; 15'h1BAB: d <= 8'hC0;
                15'h1BAC: d <= 8'hC0; 15'h1BAD: d <= 8'hC0; 15'h1BAE: d <= 8'hC0; 15'h1BAF: d <= 8'hC0;
                15'h1BB0: d <= 8'hC0; 15'h1BB1: d <= 8'hC0; 15'h1BB2: d <= 8'hC0; 15'h1BB3: d <= 8'hC0;
                15'h1BB4: d <= 8'hC0; 15'h1BB5: d <= 8'hC0; 15'h1BB6: d <= 8'hC0; 15'h1BB7: d <= 8'hC0;
                15'h1BB8: d <= 8'hC0; 15'h1BB9: d <= 8'hC0; 15'h1BBA: d <= 8'hC0; 15'h1BBB: d <= 8'hC0;
                15'h1BBC: d <= 8'hC0; 15'h1BBD: d <= 8'hC0; 15'h1BBE: d <= 8'hC0; 15'h1BBF: d <= 8'hC0;
                15'h1BC0: d <= 8'hC0; 15'h1BC1: d <= 8'hC0; 15'h1BC2: d <= 8'hC0; 15'h1BC3: d <= 8'hC0;
                15'h1BC4: d <= 8'hC0; 15'h1BC5: d <= 8'hC0; 15'h1BC6: d <= 8'hC0; 15'h1BC7: d <= 8'hC0;
                15'h1BC8: d <= 8'hC0; 15'h1BC9: d <= 8'hC0; 15'h1BCA: d <= 8'hC0; 15'h1BCB: d <= 8'hC0;
                15'h1BCC: d <= 8'hC0; 15'h1BCD: d <= 8'hC0; 15'h1BCE: d <= 8'hC0; 15'h1BCF: d <= 8'hC0;
                15'h1BD0: d <= 8'hC0; 15'h1BD1: d <= 8'hC0; 15'h1BD2: d <= 8'hC0; 15'h1BD3: d <= 8'hC0;
                15'h1BD4: d <= 8'hC0; 15'h1BD5: d <= 8'hC0; 15'h1BD6: d <= 8'hC0; 15'h1BD7: d <= 8'hC0;
                15'h1BD8: d <= 8'hC0; 15'h1BD9: d <= 8'hC0; 15'h1BDA: d <= 8'hC0; 15'h1BDB: d <= 8'hC0;
                15'h1BDC: d <= 8'hC0; 15'h1BDD: d <= 8'hC0; 15'h1BDE: d <= 8'hC0; 15'h1BDF: d <= 8'hC0;
                15'h1BE0: d <= 8'hC0; 15'h1BE1: d <= 8'hC0; 15'h1BE2: d <= 8'hC0; 15'h1BE3: d <= 8'hC0;
                15'h1BE4: d <= 8'hC0; 15'h1BE5: d <= 8'hC0; 15'h1BE6: d <= 8'hC0; 15'h1BE7: d <= 8'hC0;
                15'h1BE8: d <= 8'hC0; 15'h1BE9: d <= 8'hC0; 15'h1BEA: d <= 8'hC0; 15'h1BEB: d <= 8'hC0;
                15'h1BEC: d <= 8'hC0; 15'h1BED: d <= 8'hC0; 15'h1BEE: d <= 8'hC0; 15'h1BEF: d <= 8'hC0;
                15'h1BF0: d <= 8'hC0; 15'h1BF1: d <= 8'hC0; 15'h1BF2: d <= 8'hC0; 15'h1BF3: d <= 8'hC0;
                15'h1BF4: d <= 8'hC0; 15'h1BF5: d <= 8'hC0; 15'h1BF6: d <= 8'hC0; 15'h1BF7: d <= 8'hC0;
                15'h1BF8: d <= 8'hC0; 15'h1BF9: d <= 8'hC0; 15'h1BFA: d <= 8'hC0; 15'h1BFB: d <= 8'hC0;
                15'h1BFC: d <= 8'hC0; 15'h1BFD: d <= 8'hC0; 15'h1BFE: d <= 8'hC0; 15'h1BFF: d <= 8'hC0;
                15'h1C00: d <= 8'hC0; 15'h1C01: d <= 8'hC0; 15'h1C02: d <= 8'hC0; 15'h1C03: d <= 8'hC0;
                15'h1C04: d <= 8'hC0; 15'h1C05: d <= 8'hC0; 15'h1C06: d <= 8'hC0; 15'h1C07: d <= 8'hC0;
                15'h1C08: d <= 8'hC0; 15'h1C09: d <= 8'hC0; 15'h1C0A: d <= 8'hC0; 15'h1C0B: d <= 8'hC0;
                15'h1C0C: d <= 8'hC0; 15'h1C0D: d <= 8'hC0; 15'h1C0E: d <= 8'hC0; 15'h1C0F: d <= 8'hC0;
                15'h1C10: d <= 8'hC0; 15'h1C11: d <= 8'hC0; 15'h1C12: d <= 8'hC0; 15'h1C13: d <= 8'hC0;
                15'h1C14: d <= 8'hC0; 15'h1C15: d <= 8'hC0; 15'h1C16: d <= 8'hC0; 15'h1C17: d <= 8'hC0;
                15'h1C18: d <= 8'hC0; 15'h1C19: d <= 8'hC0; 15'h1C1A: d <= 8'hC0; 15'h1C1B: d <= 8'hC0;
                15'h1C1C: d <= 8'hC0; 15'h1C1D: d <= 8'hC0; 15'h1C1E: d <= 8'hC0; 15'h1C1F: d <= 8'hC0;
                15'h1C20: d <= 8'hC0; 15'h1C21: d <= 8'hC0; 15'h1C22: d <= 8'hC0; 15'h1C23: d <= 8'hC0;
                15'h1C24: d <= 8'hC0; 15'h1C25: d <= 8'hC0; 15'h1C26: d <= 8'hC0; 15'h1C27: d <= 8'hC0;
                15'h1C28: d <= 8'hC0; 15'h1C29: d <= 8'hC0; 15'h1C2A: d <= 8'hC0; 15'h1C2B: d <= 8'hC0;
                15'h1C2C: d <= 8'hC0; 15'h1C2D: d <= 8'hC0; 15'h1C2E: d <= 8'hC0; 15'h1C2F: d <= 8'hC0;
                15'h1C30: d <= 8'hC0; 15'h1C31: d <= 8'hC0; 15'h1C32: d <= 8'hC0; 15'h1C33: d <= 8'hC0;
                15'h1C34: d <= 8'hC0; 15'h1C35: d <= 8'hC0; 15'h1C36: d <= 8'hC0; 15'h1C37: d <= 8'hC0;
                15'h1C38: d <= 8'hC0; 15'h1C39: d <= 8'hC0; 15'h1C3A: d <= 8'hC0; 15'h1C3B: d <= 8'hC0;
                15'h1C3C: d <= 8'hC0; 15'h1C3D: d <= 8'hC0; 15'h1C3E: d <= 8'hC0; 15'h1C3F: d <= 8'hC0;
                15'h1C40: d <= 8'hC0; 15'h1C41: d <= 8'hC0; 15'h1C42: d <= 8'hC0; 15'h1C43: d <= 8'hC0;
                15'h1C44: d <= 8'hC0; 15'h1C45: d <= 8'hC0; 15'h1C46: d <= 8'hC0; 15'h1C47: d <= 8'hC0;
                15'h1C48: d <= 8'hC0; 15'h1C49: d <= 8'hC0; 15'h1C4A: d <= 8'hC0; 15'h1C4B: d <= 8'hC0;
                15'h1C4C: d <= 8'hC0; 15'h1C4D: d <= 8'hC0; 15'h1C4E: d <= 8'hC0; 15'h1C4F: d <= 8'hC0;
                15'h1C50: d <= 8'hC0; 15'h1C51: d <= 8'hC0; 15'h1C52: d <= 8'hC0; 15'h1C53: d <= 8'hC0;
                15'h1C54: d <= 8'hC0; 15'h1C55: d <= 8'hC0; 15'h1C56: d <= 8'hC0; 15'h1C57: d <= 8'hC0;
                15'h1C58: d <= 8'hC0; 15'h1C59: d <= 8'hC0; 15'h1C5A: d <= 8'hC0; 15'h1C5B: d <= 8'hC0;
                15'h1C5C: d <= 8'hC0; 15'h1C5D: d <= 8'hC0; 15'h1C5E: d <= 8'hC0; 15'h1C5F: d <= 8'hC0;
                15'h1C60: d <= 8'hC0; 15'h1C61: d <= 8'hC0; 15'h1C62: d <= 8'hC0; 15'h1C63: d <= 8'hC0;
                15'h1C64: d <= 8'hC0; 15'h1C65: d <= 8'hC0; 15'h1C66: d <= 8'hC0; 15'h1C67: d <= 8'hC0;
                15'h1C68: d <= 8'hC0; 15'h1C69: d <= 8'hC0; 15'h1C6A: d <= 8'hC0; 15'h1C6B: d <= 8'hC0;
                15'h1C6C: d <= 8'hC0; 15'h1C6D: d <= 8'hC0; 15'h1C6E: d <= 8'hC0; 15'h1C6F: d <= 8'hC0;
                15'h1C70: d <= 8'hC0; 15'h1C71: d <= 8'hC0; 15'h1C72: d <= 8'hC0; 15'h1C73: d <= 8'hC0;
                15'h1C74: d <= 8'hC0; 15'h1C75: d <= 8'hC0; 15'h1C76: d <= 8'hC0; 15'h1C77: d <= 8'hC0;
                15'h1C78: d <= 8'hC0; 15'h1C79: d <= 8'hC0; 15'h1C7A: d <= 8'hC0; 15'h1C7B: d <= 8'hC0;
                15'h1C7C: d <= 8'hC0; 15'h1C7D: d <= 8'hC0; 15'h1C7E: d <= 8'hC0; 15'h1C7F: d <= 8'hC0;
                15'h1C80: d <= 8'hC0; 15'h1C81: d <= 8'hC0; 15'h1C82: d <= 8'hC0; 15'h1C83: d <= 8'hC0;
                15'h1C84: d <= 8'hC0; 15'h1C85: d <= 8'hC0; 15'h1C86: d <= 8'hC0; 15'h1C87: d <= 8'hC0;
                15'h1C88: d <= 8'hC0; 15'h1C89: d <= 8'hC0; 15'h1C8A: d <= 8'hC0; 15'h1C8B: d <= 8'hC0;
                15'h1C8C: d <= 8'hC0; 15'h1C8D: d <= 8'hC0; 15'h1C8E: d <= 8'hC0; 15'h1C8F: d <= 8'hC0;
                15'h1C90: d <= 8'hC0; 15'h1C91: d <= 8'hC0; 15'h1C92: d <= 8'hC0; 15'h1C93: d <= 8'hC0;
                15'h1C94: d <= 8'hC0; 15'h1C95: d <= 8'hC0; 15'h1C96: d <= 8'hC0; 15'h1C97: d <= 8'hC0;
                15'h1C98: d <= 8'hC0; 15'h1C99: d <= 8'hC0; 15'h1C9A: d <= 8'hC0; 15'h1C9B: d <= 8'hC0;
                15'h1C9C: d <= 8'hC0; 15'h1C9D: d <= 8'hC0; 15'h1C9E: d <= 8'hC0; 15'h1C9F: d <= 8'hC0;
                15'h1CA0: d <= 8'hC0; 15'h1CA1: d <= 8'hC0; 15'h1CA2: d <= 8'hC0; 15'h1CA3: d <= 8'hC0;
                15'h1CA4: d <= 8'hC0; 15'h1CA5: d <= 8'hC0; 15'h1CA6: d <= 8'hC0; 15'h1CA7: d <= 8'hC0;
                15'h1CA8: d <= 8'hC0; 15'h1CA9: d <= 8'hC0; 15'h1CAA: d <= 8'hC0; 15'h1CAB: d <= 8'hC0;
                15'h1CAC: d <= 8'hC0; 15'h1CAD: d <= 8'hC0; 15'h1CAE: d <= 8'hC0; 15'h1CAF: d <= 8'hC0;
                15'h1CB0: d <= 8'hC0; 15'h1CB1: d <= 8'hC0; 15'h1CB2: d <= 8'hC0; 15'h1CB3: d <= 8'hC0;
                15'h1CB4: d <= 8'hC0; 15'h1CB5: d <= 8'hC0; 15'h1CB6: d <= 8'hC0; 15'h1CB7: d <= 8'hC0;
                15'h1CB8: d <= 8'hC0; 15'h1CB9: d <= 8'hC0; 15'h1CBA: d <= 8'hC0; 15'h1CBB: d <= 8'hC0;
                15'h1CBC: d <= 8'hC0; 15'h1CBD: d <= 8'hC0; 15'h1CBE: d <= 8'hC0; 15'h1CBF: d <= 8'hC0;
                15'h1CC0: d <= 8'hC0; 15'h1CC1: d <= 8'hC0; 15'h1CC2: d <= 8'hC0; 15'h1CC3: d <= 8'hC0;
                15'h1CC4: d <= 8'hC0; 15'h1CC5: d <= 8'hC0; 15'h1CC6: d <= 8'hC0; 15'h1CC7: d <= 8'hC0;
                15'h1CC8: d <= 8'hC0; 15'h1CC9: d <= 8'hC0; 15'h1CCA: d <= 8'hC0; 15'h1CCB: d <= 8'hC0;
                15'h1CCC: d <= 8'hC0; 15'h1CCD: d <= 8'hC0; 15'h1CCE: d <= 8'hC0; 15'h1CCF: d <= 8'hC0;
                15'h1CD0: d <= 8'hC0; 15'h1CD1: d <= 8'hC0; 15'h1CD2: d <= 8'hC0; 15'h1CD3: d <= 8'hC0;
                15'h1CD4: d <= 8'hC0; 15'h1CD5: d <= 8'hC0; 15'h1CD6: d <= 8'hC0; 15'h1CD7: d <= 8'hC0;
                15'h1CD8: d <= 8'hC0; 15'h1CD9: d <= 8'hC0; 15'h1CDA: d <= 8'hC0; 15'h1CDB: d <= 8'hC0;
                15'h1CDC: d <= 8'hC0; 15'h1CDD: d <= 8'hC0; 15'h1CDE: d <= 8'hC0; 15'h1CDF: d <= 8'hC0;
                15'h1CE0: d <= 8'hC0; 15'h1CE1: d <= 8'hC0; 15'h1CE2: d <= 8'hC0; 15'h1CE3: d <= 8'hC0;
                15'h1CE4: d <= 8'hC0; 15'h1CE5: d <= 8'hC0; 15'h1CE6: d <= 8'hC0; 15'h1CE7: d <= 8'hC0;
                15'h1CE8: d <= 8'hC0; 15'h1CE9: d <= 8'hC0; 15'h1CEA: d <= 8'hC0; 15'h1CEB: d <= 8'hC0;
                15'h1CEC: d <= 8'hC0; 15'h1CED: d <= 8'hC0; 15'h1CEE: d <= 8'hC0; 15'h1CEF: d <= 8'hC0;
                15'h1CF0: d <= 8'hC0; 15'h1CF1: d <= 8'hC0; 15'h1CF2: d <= 8'hC0; 15'h1CF3: d <= 8'hC0;
                15'h1CF4: d <= 8'hC0; 15'h1CF5: d <= 8'hC0; 15'h1CF6: d <= 8'hC0; 15'h1CF7: d <= 8'hC0;
                15'h1CF8: d <= 8'hC0; 15'h1CF9: d <= 8'hC0; 15'h1CFA: d <= 8'hC0; 15'h1CFB: d <= 8'hC0;
                15'h1CFC: d <= 8'hC0; 15'h1CFD: d <= 8'hC0; 15'h1CFE: d <= 8'hC0; 15'h1CFF: d <= 8'hC0;
                15'h1D00: d <= 8'hC0; 15'h1D01: d <= 8'hC0; 15'h1D02: d <= 8'hC0; 15'h1D03: d <= 8'hC0;
                15'h1D04: d <= 8'hC0; 15'h1D05: d <= 8'hC0; 15'h1D06: d <= 8'hC0; 15'h1D07: d <= 8'hC0;
                15'h1D08: d <= 8'hC0; 15'h1D09: d <= 8'hC0; 15'h1D0A: d <= 8'hC0; 15'h1D0B: d <= 8'hC0;
                15'h1D0C: d <= 8'hC0; 15'h1D0D: d <= 8'hC0; 15'h1D0E: d <= 8'hC0; 15'h1D0F: d <= 8'hC0;
                15'h1D10: d <= 8'hC0; 15'h1D11: d <= 8'hC0; 15'h1D12: d <= 8'hC0; 15'h1D13: d <= 8'hC0;
                15'h1D14: d <= 8'hC0; 15'h1D15: d <= 8'hC0; 15'h1D16: d <= 8'hC0; 15'h1D17: d <= 8'hC0;
                15'h1D18: d <= 8'hC0; 15'h1D19: d <= 8'hC0; 15'h1D1A: d <= 8'hC0; 15'h1D1B: d <= 8'hC0;
                15'h1D1C: d <= 8'hC0; 15'h1D1D: d <= 8'hC0; 15'h1D1E: d <= 8'hC0; 15'h1D1F: d <= 8'hC0;
                15'h1D20: d <= 8'hC0; 15'h1D21: d <= 8'hC0; 15'h1D22: d <= 8'hC0; 15'h1D23: d <= 8'hC0;
                15'h1D24: d <= 8'hC0; 15'h1D25: d <= 8'hC0; 15'h1D26: d <= 8'hC0; 15'h1D27: d <= 8'hC0;
                15'h1D28: d <= 8'hC0; 15'h1D29: d <= 8'hC0; 15'h1D2A: d <= 8'hC0; 15'h1D2B: d <= 8'hC0;
                15'h1D2C: d <= 8'hC0; 15'h1D2D: d <= 8'hC0; 15'h1D2E: d <= 8'hC0; 15'h1D2F: d <= 8'hC0;
                15'h1D30: d <= 8'hC0; 15'h1D31: d <= 8'hC0; 15'h1D32: d <= 8'hC0; 15'h1D33: d <= 8'hC0;
                15'h1D34: d <= 8'hC0; 15'h1D35: d <= 8'hC0; 15'h1D36: d <= 8'hC0; 15'h1D37: d <= 8'hC0;
                15'h1D38: d <= 8'hC0; 15'h1D39: d <= 8'hC0; 15'h1D3A: d <= 8'hC0; 15'h1D3B: d <= 8'hC0;
                15'h1D3C: d <= 8'hC0; 15'h1D3D: d <= 8'hC0; 15'h1D3E: d <= 8'hC0; 15'h1D3F: d <= 8'hC0;
                15'h1D40: d <= 8'hC0; 15'h1D41: d <= 8'hC0; 15'h1D42: d <= 8'hC0; 15'h1D43: d <= 8'hC0;
                15'h1D44: d <= 8'hC0; 15'h1D45: d <= 8'hC0; 15'h1D46: d <= 8'hC0; 15'h1D47: d <= 8'hC0;
                15'h1D48: d <= 8'hC0; 15'h1D49: d <= 8'hC0; 15'h1D4A: d <= 8'hC0; 15'h1D4B: d <= 8'hC0;
                15'h1D4C: d <= 8'hC0; 15'h1D4D: d <= 8'hC0; 15'h1D4E: d <= 8'hC0; 15'h1D4F: d <= 8'hC0;
                15'h1D50: d <= 8'hC0; 15'h1D51: d <= 8'hC0; 15'h1D52: d <= 8'hC0; 15'h1D53: d <= 8'hC0;
                15'h1D54: d <= 8'hC0; 15'h1D55: d <= 8'hC0; 15'h1D56: d <= 8'hC0; 15'h1D57: d <= 8'hC0;
                15'h1D58: d <= 8'hC0; 15'h1D59: d <= 8'hC0; 15'h1D5A: d <= 8'hC0; 15'h1D5B: d <= 8'hC0;
                15'h1D5C: d <= 8'hC0; 15'h1D5D: d <= 8'hC0; 15'h1D5E: d <= 8'hC0; 15'h1D5F: d <= 8'hC0;
                15'h1D60: d <= 8'hC0; 15'h1D61: d <= 8'hC0; 15'h1D62: d <= 8'hC0; 15'h1D63: d <= 8'hC0;
                15'h1D64: d <= 8'hC0; 15'h1D65: d <= 8'hC0; 15'h1D66: d <= 8'hC0; 15'h1D67: d <= 8'hC0;
                15'h1D68: d <= 8'hC0; 15'h1D69: d <= 8'hC0; 15'h1D6A: d <= 8'hC0; 15'h1D6B: d <= 8'hC0;
                15'h1D6C: d <= 8'hC0; 15'h1D6D: d <= 8'hC0; 15'h1D6E: d <= 8'hC0; 15'h1D6F: d <= 8'hC0;
                15'h1D70: d <= 8'hC0; 15'h1D71: d <= 8'hC0; 15'h1D72: d <= 8'hC0; 15'h1D73: d <= 8'hC0;
                15'h1D74: d <= 8'hC0; 15'h1D75: d <= 8'hC0; 15'h1D76: d <= 8'hC0; 15'h1D77: d <= 8'hC0;
                15'h1D78: d <= 8'hC0; 15'h1D79: d <= 8'hC0; 15'h1D7A: d <= 8'hC0; 15'h1D7B: d <= 8'hC0;
                15'h1D7C: d <= 8'hC0; 15'h1D7D: d <= 8'hC0; 15'h1D7E: d <= 8'hC0; 15'h1D7F: d <= 8'hC0;
                15'h1D80: d <= 8'hC0; 15'h1D81: d <= 8'hC0; 15'h1D82: d <= 8'hC0; 15'h1D83: d <= 8'hC0;
                15'h1D84: d <= 8'hC0; 15'h1D85: d <= 8'hC0; 15'h1D86: d <= 8'hC0; 15'h1D87: d <= 8'hC0;
                15'h1D88: d <= 8'hC0; 15'h1D89: d <= 8'hC0; 15'h1D8A: d <= 8'hC0; 15'h1D8B: d <= 8'hC0;
                15'h1D8C: d <= 8'hC0; 15'h1D8D: d <= 8'hC0; 15'h1D8E: d <= 8'hC0; 15'h1D8F: d <= 8'hC0;
                15'h1D90: d <= 8'hC0; 15'h1D91: d <= 8'hC0; 15'h1D92: d <= 8'hC0; 15'h1D93: d <= 8'hC0;
                15'h1D94: d <= 8'hC0; 15'h1D95: d <= 8'hC0; 15'h1D96: d <= 8'hC0; 15'h1D97: d <= 8'hC0;
                15'h1D98: d <= 8'hC0; 15'h1D99: d <= 8'hC0; 15'h1D9A: d <= 8'hC0; 15'h1D9B: d <= 8'hC0;
                15'h1D9C: d <= 8'hC0; 15'h1D9D: d <= 8'hC0; 15'h1D9E: d <= 8'hC0; 15'h1D9F: d <= 8'hC0;
                15'h1DA0: d <= 8'hC0; 15'h1DA1: d <= 8'hC0; 15'h1DA2: d <= 8'hC0; 15'h1DA3: d <= 8'hC0;
                15'h1DA4: d <= 8'hC0; 15'h1DA5: d <= 8'hC0; 15'h1DA6: d <= 8'hC0; 15'h1DA7: d <= 8'hC0;
                15'h1DA8: d <= 8'hC0; 15'h1DA9: d <= 8'hC0; 15'h1DAA: d <= 8'hC0; 15'h1DAB: d <= 8'hC0;
                15'h1DAC: d <= 8'hC0; 15'h1DAD: d <= 8'hC0; 15'h1DAE: d <= 8'hC0; 15'h1DAF: d <= 8'hC0;
                15'h1DB0: d <= 8'hC0; 15'h1DB1: d <= 8'hC0; 15'h1DB2: d <= 8'hC0; 15'h1DB3: d <= 8'hC0;
                15'h1DB4: d <= 8'hC0; 15'h1DB5: d <= 8'hC0; 15'h1DB6: d <= 8'hC0; 15'h1DB7: d <= 8'hC0;
                15'h1DB8: d <= 8'hC0; 15'h1DB9: d <= 8'hC0; 15'h1DBA: d <= 8'hC0; 15'h1DBB: d <= 8'hC0;
                15'h1DBC: d <= 8'hC0; 15'h1DBD: d <= 8'hC0; 15'h1DBE: d <= 8'hC0; 15'h1DBF: d <= 8'hC0;
                15'h1DC0: d <= 8'hC0; 15'h1DC1: d <= 8'hC0; 15'h1DC2: d <= 8'hC0; 15'h1DC3: d <= 8'hC0;
                15'h1DC4: d <= 8'hC0; 15'h1DC5: d <= 8'hC0; 15'h1DC6: d <= 8'hC0; 15'h1DC7: d <= 8'hC0;
                15'h1DC8: d <= 8'hC0; 15'h1DC9: d <= 8'hC0; 15'h1DCA: d <= 8'hC0; 15'h1DCB: d <= 8'hC0;
                15'h1DCC: d <= 8'hC0; 15'h1DCD: d <= 8'hC0; 15'h1DCE: d <= 8'hC0; 15'h1DCF: d <= 8'hC0;
                15'h1DD0: d <= 8'hC0; 15'h1DD1: d <= 8'hC0; 15'h1DD2: d <= 8'hC0; 15'h1DD3: d <= 8'hC0;
                15'h1DD4: d <= 8'hC0; 15'h1DD5: d <= 8'hC0; 15'h1DD6: d <= 8'hC0; 15'h1DD7: d <= 8'hC0;
                15'h1DD8: d <= 8'hC0; 15'h1DD9: d <= 8'hC0; 15'h1DDA: d <= 8'hC0; 15'h1DDB: d <= 8'hC0;
                15'h1DDC: d <= 8'hC0; 15'h1DDD: d <= 8'hC0; 15'h1DDE: d <= 8'hC0; 15'h1DDF: d <= 8'hC0;
                15'h1DE0: d <= 8'hC0; 15'h1DE1: d <= 8'hC0; 15'h1DE2: d <= 8'hC0; 15'h1DE3: d <= 8'hC0;
                15'h1DE4: d <= 8'hC0; 15'h1DE5: d <= 8'hC0; 15'h1DE6: d <= 8'hC0; 15'h1DE7: d <= 8'hC0;
                15'h1DE8: d <= 8'hC0; 15'h1DE9: d <= 8'hC0; 15'h1DEA: d <= 8'hC0; 15'h1DEB: d <= 8'hC0;
                15'h1DEC: d <= 8'hC0; 15'h1DED: d <= 8'hC0; 15'h1DEE: d <= 8'hC0; 15'h1DEF: d <= 8'hC0;
                15'h1DF0: d <= 8'hC0; 15'h1DF1: d <= 8'hC0; 15'h1DF2: d <= 8'hC0; 15'h1DF3: d <= 8'hC0;
                15'h1DF4: d <= 8'hC0; 15'h1DF5: d <= 8'hC0; 15'h1DF6: d <= 8'hC0; 15'h1DF7: d <= 8'hC0;
                15'h1DF8: d <= 8'hC0; 15'h1DF9: d <= 8'hC0; 15'h1DFA: d <= 8'hC0; 15'h1DFB: d <= 8'hC0;
                15'h1DFC: d <= 8'hC0; 15'h1DFD: d <= 8'hC0; 15'h1DFE: d <= 8'hC0; 15'h1DFF: d <= 8'hC0;
                15'h1E00: d <= 8'hC0; 15'h1E01: d <= 8'hC0; 15'h1E02: d <= 8'hC0; 15'h1E03: d <= 8'hC0;
                15'h1E04: d <= 8'hC0; 15'h1E05: d <= 8'hC0; 15'h1E06: d <= 8'hC0; 15'h1E07: d <= 8'hC0;
                15'h1E08: d <= 8'hC0; 15'h1E09: d <= 8'hC0; 15'h1E0A: d <= 8'hC0; 15'h1E0B: d <= 8'hC0;
                15'h1E0C: d <= 8'hC0; 15'h1E0D: d <= 8'hC0; 15'h1E0E: d <= 8'hC0; 15'h1E0F: d <= 8'hC0;
                15'h1E10: d <= 8'hC0; 15'h1E11: d <= 8'hC0; 15'h1E12: d <= 8'hC0; 15'h1E13: d <= 8'hC0;
                15'h1E14: d <= 8'hC0; 15'h1E15: d <= 8'hC0; 15'h1E16: d <= 8'hC0; 15'h1E17: d <= 8'hC0;
                15'h1E18: d <= 8'hC0; 15'h1E19: d <= 8'hC0; 15'h1E1A: d <= 8'hC0; 15'h1E1B: d <= 8'hC0;
                15'h1E1C: d <= 8'hC0; 15'h1E1D: d <= 8'hC0; 15'h1E1E: d <= 8'hC0; 15'h1E1F: d <= 8'hC0;
                15'h1E20: d <= 8'hC0; 15'h1E21: d <= 8'hC0; 15'h1E22: d <= 8'hC0; 15'h1E23: d <= 8'hC0;
                15'h1E24: d <= 8'hC0; 15'h1E25: d <= 8'hC0; 15'h1E26: d <= 8'hC0; 15'h1E27: d <= 8'hC0;
                15'h1E28: d <= 8'hC0; 15'h1E29: d <= 8'hC0; 15'h1E2A: d <= 8'hC0; 15'h1E2B: d <= 8'hC0;
                15'h1E2C: d <= 8'hC0; 15'h1E2D: d <= 8'hC0; 15'h1E2E: d <= 8'hC0; 15'h1E2F: d <= 8'hC0;
                15'h1E30: d <= 8'hC0; 15'h1E31: d <= 8'hC0; 15'h1E32: d <= 8'hC0; 15'h1E33: d <= 8'hC0;
                15'h1E34: d <= 8'hC0; 15'h1E35: d <= 8'hC0; 15'h1E36: d <= 8'hC0; 15'h1E37: d <= 8'hC0;
                15'h1E38: d <= 8'hC0; 15'h1E39: d <= 8'hC0; 15'h1E3A: d <= 8'hC0; 15'h1E3B: d <= 8'hC0;
                15'h1E3C: d <= 8'hC0; 15'h1E3D: d <= 8'hC0; 15'h1E3E: d <= 8'hC0; 15'h1E3F: d <= 8'hC0;
                15'h1E40: d <= 8'hC0; 15'h1E41: d <= 8'hC0; 15'h1E42: d <= 8'hC0; 15'h1E43: d <= 8'hC0;
                15'h1E44: d <= 8'hC0; 15'h1E45: d <= 8'hC0; 15'h1E46: d <= 8'hC0; 15'h1E47: d <= 8'hC0;
                15'h1E48: d <= 8'hC0; 15'h1E49: d <= 8'hC0; 15'h1E4A: d <= 8'hC0; 15'h1E4B: d <= 8'hC0;
                15'h1E4C: d <= 8'hC0; 15'h1E4D: d <= 8'hC0; 15'h1E4E: d <= 8'hC0; 15'h1E4F: d <= 8'hC0;
                15'h1E50: d <= 8'hC0; 15'h1E51: d <= 8'hC0; 15'h1E52: d <= 8'hC0; 15'h1E53: d <= 8'hC0;
                15'h1E54: d <= 8'hC0; 15'h1E55: d <= 8'hC0; 15'h1E56: d <= 8'hC0; 15'h1E57: d <= 8'hC0;
                15'h1E58: d <= 8'hC0; 15'h1E59: d <= 8'hC0; 15'h1E5A: d <= 8'hC0; 15'h1E5B: d <= 8'hC0;
                15'h1E5C: d <= 8'hC0; 15'h1E5D: d <= 8'hC0; 15'h1E5E: d <= 8'hC0; 15'h1E5F: d <= 8'hC0;
                15'h1E60: d <= 8'hC0; 15'h1E61: d <= 8'hC0; 15'h1E62: d <= 8'hC0; 15'h1E63: d <= 8'hC0;
                15'h1E64: d <= 8'hC0; 15'h1E65: d <= 8'hC0; 15'h1E66: d <= 8'hC0; 15'h1E67: d <= 8'hC0;
                15'h1E68: d <= 8'hC0; 15'h1E69: d <= 8'hC0; 15'h1E6A: d <= 8'hC0; 15'h1E6B: d <= 8'hC0;
                15'h1E6C: d <= 8'hC0; 15'h1E6D: d <= 8'hC0; 15'h1E6E: d <= 8'hC0; 15'h1E6F: d <= 8'hC0;
                15'h1E70: d <= 8'hC0; 15'h1E71: d <= 8'hC0; 15'h1E72: d <= 8'hC0; 15'h1E73: d <= 8'hC0;
                15'h1E74: d <= 8'hC0; 15'h1E75: d <= 8'hC0; 15'h1E76: d <= 8'hC0; 15'h1E77: d <= 8'hC0;
                15'h1E78: d <= 8'hC0; 15'h1E79: d <= 8'hC0; 15'h1E7A: d <= 8'hC0; 15'h1E7B: d <= 8'hC0;
                15'h1E7C: d <= 8'hC0; 15'h1E7D: d <= 8'hC0; 15'h1E7E: d <= 8'hC0; 15'h1E7F: d <= 8'hC0;
                15'h1E80: d <= 8'hC0; 15'h1E81: d <= 8'hC0; 15'h1E82: d <= 8'hC0; 15'h1E83: d <= 8'hC0;
                15'h1E84: d <= 8'hC0; 15'h1E85: d <= 8'hC0; 15'h1E86: d <= 8'hC0; 15'h1E87: d <= 8'hC0;
                15'h1E88: d <= 8'hC0; 15'h1E89: d <= 8'hC0; 15'h1E8A: d <= 8'hC0; 15'h1E8B: d <= 8'hC0;
                15'h1E8C: d <= 8'hC0; 15'h1E8D: d <= 8'hC0; 15'h1E8E: d <= 8'hC0; 15'h1E8F: d <= 8'hC0;
                15'h1E90: d <= 8'hC0; 15'h1E91: d <= 8'hC0; 15'h1E92: d <= 8'hC0; 15'h1E93: d <= 8'hC0;
                15'h1E94: d <= 8'hC0; 15'h1E95: d <= 8'hC0; 15'h1E96: d <= 8'hC0; 15'h1E97: d <= 8'hC0;
                15'h1E98: d <= 8'hC0; 15'h1E99: d <= 8'hC0; 15'h1E9A: d <= 8'hC0; 15'h1E9B: d <= 8'hC0;
                15'h1E9C: d <= 8'hC0; 15'h1E9D: d <= 8'hC0; 15'h1E9E: d <= 8'hC0; 15'h1E9F: d <= 8'hC0;
                15'h1EA0: d <= 8'hC0; 15'h1EA1: d <= 8'hC0; 15'h1EA2: d <= 8'hC0; 15'h1EA3: d <= 8'hC0;
                15'h1EA4: d <= 8'hC0; 15'h1EA5: d <= 8'hC0; 15'h1EA6: d <= 8'hC0; 15'h1EA7: d <= 8'hC0;
                15'h1EA8: d <= 8'hC0; 15'h1EA9: d <= 8'hC0; 15'h1EAA: d <= 8'hC0; 15'h1EAB: d <= 8'hC0;
                15'h1EAC: d <= 8'hC0; 15'h1EAD: d <= 8'hC0; 15'h1EAE: d <= 8'hC0; 15'h1EAF: d <= 8'hC0;
                15'h1EB0: d <= 8'hC0; 15'h1EB1: d <= 8'hC0; 15'h1EB2: d <= 8'hC0; 15'h1EB3: d <= 8'hC0;
                15'h1EB4: d <= 8'hC0; 15'h1EB5: d <= 8'hC0; 15'h1EB6: d <= 8'hC0; 15'h1EB7: d <= 8'hC0;
                15'h1EB8: d <= 8'hC0; 15'h1EB9: d <= 8'hC0; 15'h1EBA: d <= 8'hC0; 15'h1EBB: d <= 8'hC0;
                15'h1EBC: d <= 8'hC0; 15'h1EBD: d <= 8'hC0; 15'h1EBE: d <= 8'hC0; 15'h1EBF: d <= 8'hC0;
                15'h1EC0: d <= 8'hC0; 15'h1EC1: d <= 8'hC0; 15'h1EC2: d <= 8'hC0; 15'h1EC3: d <= 8'hC0;
                15'h1EC4: d <= 8'hC0; 15'h1EC5: d <= 8'hC0; 15'h1EC6: d <= 8'hC0; 15'h1EC7: d <= 8'hC0;
                15'h1EC8: d <= 8'hC0; 15'h1EC9: d <= 8'hC0; 15'h1ECA: d <= 8'hC0; 15'h1ECB: d <= 8'hC0;
                15'h1ECC: d <= 8'hC0; 15'h1ECD: d <= 8'hC0; 15'h1ECE: d <= 8'hC0; 15'h1ECF: d <= 8'hC0;
                15'h1ED0: d <= 8'hC0; 15'h1ED1: d <= 8'hC0; 15'h1ED2: d <= 8'hC0; 15'h1ED3: d <= 8'hC0;
                15'h1ED4: d <= 8'hC0; 15'h1ED5: d <= 8'hC0; 15'h1ED6: d <= 8'hC0; 15'h1ED7: d <= 8'hC0;
                15'h1ED8: d <= 8'hC0; 15'h1ED9: d <= 8'hC0; 15'h1EDA: d <= 8'hC0; 15'h1EDB: d <= 8'hC0;
                15'h1EDC: d <= 8'hC0; 15'h1EDD: d <= 8'hC0; 15'h1EDE: d <= 8'hC0; 15'h1EDF: d <= 8'hC0;
                15'h1EE0: d <= 8'hC0; 15'h1EE1: d <= 8'hC0; 15'h1EE2: d <= 8'hC0; 15'h1EE3: d <= 8'hC0;
                15'h1EE4: d <= 8'hC0; 15'h1EE5: d <= 8'hC0; 15'h1EE6: d <= 8'hC0; 15'h1EE7: d <= 8'hC0;
                15'h1EE8: d <= 8'hC0; 15'h1EE9: d <= 8'hC0; 15'h1EEA: d <= 8'hC0; 15'h1EEB: d <= 8'hC0;
                15'h1EEC: d <= 8'hC0; 15'h1EED: d <= 8'hC0; 15'h1EEE: d <= 8'hC0; 15'h1EEF: d <= 8'hC0;
                15'h1EF0: d <= 8'hC0; 15'h1EF1: d <= 8'hC0; 15'h1EF2: d <= 8'hC0; 15'h1EF3: d <= 8'hC0;
                15'h1EF4: d <= 8'hC0; 15'h1EF5: d <= 8'hC0; 15'h1EF6: d <= 8'hC0; 15'h1EF7: d <= 8'hC0;
                15'h1EF8: d <= 8'hC0; 15'h1EF9: d <= 8'hC0; 15'h1EFA: d <= 8'hC0; 15'h1EFB: d <= 8'hC0;
                15'h1EFC: d <= 8'hC0; 15'h1EFD: d <= 8'hC0; 15'h1EFE: d <= 8'hC0; 15'h1EFF: d <= 8'hC0;
                15'h1F00: d <= 8'hC0; 15'h1F01: d <= 8'hC0; 15'h1F02: d <= 8'hC0; 15'h1F03: d <= 8'hC0;
                15'h1F04: d <= 8'hC0; 15'h1F05: d <= 8'hC0; 15'h1F06: d <= 8'hC0; 15'h1F07: d <= 8'hC0;
                15'h1F08: d <= 8'hC0; 15'h1F09: d <= 8'hC0; 15'h1F0A: d <= 8'hC0; 15'h1F0B: d <= 8'hC0;
                15'h1F0C: d <= 8'hC0; 15'h1F0D: d <= 8'hC0; 15'h1F0E: d <= 8'hC0; 15'h1F0F: d <= 8'hC0;
                15'h1F10: d <= 8'hC0; 15'h1F11: d <= 8'hC0; 15'h1F12: d <= 8'hC0; 15'h1F13: d <= 8'hC0;
                15'h1F14: d <= 8'hC0; 15'h1F15: d <= 8'hC0; 15'h1F16: d <= 8'hC0; 15'h1F17: d <= 8'hC0;
                15'h1F18: d <= 8'hC0; 15'h1F19: d <= 8'hC0; 15'h1F1A: d <= 8'hC0; 15'h1F1B: d <= 8'hC0;
                15'h1F1C: d <= 8'hC0; 15'h1F1D: d <= 8'hC0; 15'h1F1E: d <= 8'hC0; 15'h1F1F: d <= 8'hC0;
                15'h1F20: d <= 8'hC0; 15'h1F21: d <= 8'hC0; 15'h1F22: d <= 8'hC0; 15'h1F23: d <= 8'hC0;
                15'h1F24: d <= 8'hC0; 15'h1F25: d <= 8'hC0; 15'h1F26: d <= 8'hC0; 15'h1F27: d <= 8'hC0;
                15'h1F28: d <= 8'hC0; 15'h1F29: d <= 8'hC0; 15'h1F2A: d <= 8'hC0; 15'h1F2B: d <= 8'hC0;
                15'h1F2C: d <= 8'hC0; 15'h1F2D: d <= 8'hC0; 15'h1F2E: d <= 8'hC0; 15'h1F2F: d <= 8'hC0;
                15'h1F30: d <= 8'hC0; 15'h1F31: d <= 8'hC0; 15'h1F32: d <= 8'hC0; 15'h1F33: d <= 8'hC0;
                15'h1F34: d <= 8'hC0; 15'h1F35: d <= 8'hC0; 15'h1F36: d <= 8'hC0; 15'h1F37: d <= 8'hC0;
                15'h1F38: d <= 8'hC0; 15'h1F39: d <= 8'hC0; 15'h1F3A: d <= 8'hC0; 15'h1F3B: d <= 8'hC0;
                15'h1F3C: d <= 8'hC0; 15'h1F3D: d <= 8'hC0; 15'h1F3E: d <= 8'hC0; 15'h1F3F: d <= 8'hC0;
                15'h1F40: d <= 8'hC0; 15'h1F41: d <= 8'hC0; 15'h1F42: d <= 8'hC0; 15'h1F43: d <= 8'hC0;
                15'h1F44: d <= 8'hC0; 15'h1F45: d <= 8'hC0; 15'h1F46: d <= 8'hC0; 15'h1F47: d <= 8'hC0;
                15'h1F48: d <= 8'hC0; 15'h1F49: d <= 8'hC0; 15'h1F4A: d <= 8'hC0; 15'h1F4B: d <= 8'hC0;
                15'h1F4C: d <= 8'hC0; 15'h1F4D: d <= 8'hC0; 15'h1F4E: d <= 8'hC0; 15'h1F4F: d <= 8'hC0;
                15'h1F50: d <= 8'hC0; 15'h1F51: d <= 8'hC0; 15'h1F52: d <= 8'hC0; 15'h1F53: d <= 8'hC0;
                15'h1F54: d <= 8'hC0; 15'h1F55: d <= 8'hC0; 15'h1F56: d <= 8'hC0; 15'h1F57: d <= 8'hC0;
                15'h1F58: d <= 8'hC0; 15'h1F59: d <= 8'hC0; 15'h1F5A: d <= 8'hC0; 15'h1F5B: d <= 8'hC0;
                15'h1F5C: d <= 8'hC0; 15'h1F5D: d <= 8'hC0; 15'h1F5E: d <= 8'hC0; 15'h1F5F: d <= 8'hC0;
                15'h1F60: d <= 8'hC0; 15'h1F61: d <= 8'hC0; 15'h1F62: d <= 8'hC0; 15'h1F63: d <= 8'hC0;
                15'h1F64: d <= 8'hC0; 15'h1F65: d <= 8'hC0; 15'h1F66: d <= 8'hC0; 15'h1F67: d <= 8'hC0;
                15'h1F68: d <= 8'hC0; 15'h1F69: d <= 8'hC0; 15'h1F6A: d <= 8'hC0; 15'h1F6B: d <= 8'hC0;
                15'h1F6C: d <= 8'hC0; 15'h1F6D: d <= 8'hC0; 15'h1F6E: d <= 8'hC0; 15'h1F6F: d <= 8'hC0;
                15'h1F70: d <= 8'hC0; 15'h1F71: d <= 8'hC0; 15'h1F72: d <= 8'hC0; 15'h1F73: d <= 8'hC0;
                15'h1F74: d <= 8'hC0; 15'h1F75: d <= 8'hC0; 15'h1F76: d <= 8'hC0; 15'h1F77: d <= 8'hC0;
                15'h1F78: d <= 8'hC0; 15'h1F79: d <= 8'hC0; 15'h1F7A: d <= 8'hC0; 15'h1F7B: d <= 8'hC0;
                15'h1F7C: d <= 8'hC0; 15'h1F7D: d <= 8'hC0; 15'h1F7E: d <= 8'hC0; 15'h1F7F: d <= 8'hC0;
                15'h1F80: d <= 8'hC0; 15'h1F81: d <= 8'hC0; 15'h1F82: d <= 8'hC0; 15'h1F83: d <= 8'hC0;
                15'h1F84: d <= 8'hC0; 15'h1F85: d <= 8'hC0; 15'h1F86: d <= 8'hC0; 15'h1F87: d <= 8'hC0;
                15'h1F88: d <= 8'hC0; 15'h1F89: d <= 8'hC0; 15'h1F8A: d <= 8'hC0; 15'h1F8B: d <= 8'hC0;
                15'h1F8C: d <= 8'hC0; 15'h1F8D: d <= 8'hC0; 15'h1F8E: d <= 8'hC0; 15'h1F8F: d <= 8'hC0;
                15'h1F90: d <= 8'hC0; 15'h1F91: d <= 8'hC0; 15'h1F92: d <= 8'hC0; 15'h1F93: d <= 8'hC0;
                15'h1F94: d <= 8'hC0; 15'h1F95: d <= 8'hC0; 15'h1F96: d <= 8'hC0; 15'h1F97: d <= 8'hC0;
                15'h1F98: d <= 8'hC0; 15'h1F99: d <= 8'hC0; 15'h1F9A: d <= 8'hC0; 15'h1F9B: d <= 8'hC0;
                15'h1F9C: d <= 8'hC0; 15'h1F9D: d <= 8'hC0; 15'h1F9E: d <= 8'hC0; 15'h1F9F: d <= 8'hC0;
                15'h1FA0: d <= 8'hC0; 15'h1FA1: d <= 8'hC0; 15'h1FA2: d <= 8'hC0; 15'h1FA3: d <= 8'hC0;
                15'h1FA4: d <= 8'hC0; 15'h1FA5: d <= 8'hC0; 15'h1FA6: d <= 8'hC0; 15'h1FA7: d <= 8'hC0;
                15'h1FA8: d <= 8'hC0; 15'h1FA9: d <= 8'hC0; 15'h1FAA: d <= 8'hC0; 15'h1FAB: d <= 8'hC0;
                15'h1FAC: d <= 8'hC0; 15'h1FAD: d <= 8'hC0; 15'h1FAE: d <= 8'hC0; 15'h1FAF: d <= 8'hC0;
                15'h1FB0: d <= 8'hC0; 15'h1FB1: d <= 8'hC0; 15'h1FB2: d <= 8'hC0; 15'h1FB3: d <= 8'hC0;
                15'h1FB4: d <= 8'hC0; 15'h1FB5: d <= 8'hC0; 15'h1FB6: d <= 8'hC0; 15'h1FB7: d <= 8'hC0;
                15'h1FB8: d <= 8'hC0; 15'h1FB9: d <= 8'hC0; 15'h1FBA: d <= 8'hC0; 15'h1FBB: d <= 8'hC0;
                15'h1FBC: d <= 8'hC0; 15'h1FBD: d <= 8'hC0; 15'h1FBE: d <= 8'hC0; 15'h1FBF: d <= 8'hC0;
                15'h1FC0: d <= 8'hC0; 15'h1FC1: d <= 8'hC0; 15'h1FC2: d <= 8'hC0; 15'h1FC3: d <= 8'hC0;
                15'h1FC4: d <= 8'hC0; 15'h1FC5: d <= 8'hC0; 15'h1FC6: d <= 8'hC0; 15'h1FC7: d <= 8'hC0;
                15'h1FC8: d <= 8'hC0; 15'h1FC9: d <= 8'hC0; 15'h1FCA: d <= 8'hC0; 15'h1FCB: d <= 8'hC0;
                15'h1FCC: d <= 8'hC0; 15'h1FCD: d <= 8'hC0; 15'h1FCE: d <= 8'hC0; 15'h1FCF: d <= 8'hC0;
                15'h1FD0: d <= 8'hC0; 15'h1FD1: d <= 8'hC0; 15'h1FD2: d <= 8'hC0; 15'h1FD3: d <= 8'hC0;
                15'h1FD4: d <= 8'hC0; 15'h1FD5: d <= 8'hC0; 15'h1FD6: d <= 8'hC0; 15'h1FD7: d <= 8'hC0;
                15'h1FD8: d <= 8'hC0; 15'h1FD9: d <= 8'hC0; 15'h1FDA: d <= 8'hC0; 15'h1FDB: d <= 8'hC0;
                15'h1FDC: d <= 8'hC0; 15'h1FDD: d <= 8'hC0; 15'h1FDE: d <= 8'hC0; 15'h1FDF: d <= 8'hC0;
                15'h1FE0: d <= 8'hC0; 15'h1FE1: d <= 8'hC0; 15'h1FE2: d <= 8'hC0; 15'h1FE3: d <= 8'hC0;
                15'h1FE4: d <= 8'hC0; 15'h1FE5: d <= 8'hC0; 15'h1FE6: d <= 8'hC0; 15'h1FE7: d <= 8'hC0;
                15'h1FE8: d <= 8'hC0; 15'h1FE9: d <= 8'hC0; 15'h1FEA: d <= 8'hC0; 15'h1FEB: d <= 8'hC0;
                15'h1FEC: d <= 8'hC0; 15'h1FED: d <= 8'hC0; 15'h1FEE: d <= 8'hC0; 15'h1FEF: d <= 8'hC0;
                15'h1FF0: d <= 8'hC0; 15'h1FF1: d <= 8'hC0; 15'h1FF2: d <= 8'hC0; 15'h1FF3: d <= 8'hC0;
                15'h1FF4: d <= 8'hC0; 15'h1FF5: d <= 8'hC0; 15'h1FF6: d <= 8'hC0; 15'h1FF7: d <= 8'hC0;
                15'h1FF8: d <= 8'hC0; 15'h1FF9: d <= 8'hC0; 15'h1FFA: d <= 8'hC0; 15'h1FFB: d <= 8'hC0;
                15'h1FFC: d <= 8'hC0; 15'h1FFD: d <= 8'hC0; 15'h1FFE: d <= 8'hC0; 15'h1FFF: d <= 8'hC0;
                15'h2000: d <= 8'hC0; 15'h2001: d <= 8'hC0; 15'h2002: d <= 8'hC0; 15'h2003: d <= 8'hC0;
                15'h2004: d <= 8'hC0; 15'h2005: d <= 8'hC0; 15'h2006: d <= 8'hC0; 15'h2007: d <= 8'hC0;
                15'h2008: d <= 8'hC0; 15'h2009: d <= 8'hC0; 15'h200A: d <= 8'hC0; 15'h200B: d <= 8'hC0;
                15'h200C: d <= 8'hC0; 15'h200D: d <= 8'hC0; 15'h200E: d <= 8'hC0; 15'h200F: d <= 8'hC0;
                15'h2010: d <= 8'hC0; 15'h2011: d <= 8'hC0; 15'h2012: d <= 8'hC0; 15'h2013: d <= 8'hC0;
                15'h2014: d <= 8'hC0; 15'h2015: d <= 8'hC0; 15'h2016: d <= 8'hC0; 15'h2017: d <= 8'hC0;
                15'h2018: d <= 8'hC0; 15'h2019: d <= 8'hC0; 15'h201A: d <= 8'hC0; 15'h201B: d <= 8'hC0;
                15'h201C: d <= 8'hC0; 15'h201D: d <= 8'hC0; 15'h201E: d <= 8'hC0; 15'h201F: d <= 8'hC0;
                15'h2020: d <= 8'hC0; 15'h2021: d <= 8'hC0; 15'h2022: d <= 8'hC0; 15'h2023: d <= 8'hC0;
                15'h2024: d <= 8'hC0; 15'h2025: d <= 8'hC0; 15'h2026: d <= 8'hC0; 15'h2027: d <= 8'hC0;
                15'h2028: d <= 8'hC0; 15'h2029: d <= 8'hC0; 15'h202A: d <= 8'hC0; 15'h202B: d <= 8'hC0;
                15'h202C: d <= 8'hC0; 15'h202D: d <= 8'hC0; 15'h202E: d <= 8'hC0; 15'h202F: d <= 8'hC0;
                15'h2030: d <= 8'hC0; 15'h2031: d <= 8'hC0; 15'h2032: d <= 8'hC0; 15'h2033: d <= 8'hC0;
                15'h2034: d <= 8'hC0; 15'h2035: d <= 8'hC0; 15'h2036: d <= 8'hC0; 15'h2037: d <= 8'hC0;
                15'h2038: d <= 8'hC0; 15'h2039: d <= 8'hC0; 15'h203A: d <= 8'hC0; 15'h203B: d <= 8'hC0;
                15'h203C: d <= 8'hC0; 15'h203D: d <= 8'hC0; 15'h203E: d <= 8'hC0; 15'h203F: d <= 8'hC0;
                15'h2040: d <= 8'hC0; 15'h2041: d <= 8'hC0; 15'h2042: d <= 8'hC0; 15'h2043: d <= 8'hC0;
                15'h2044: d <= 8'hC0; 15'h2045: d <= 8'hC0; 15'h2046: d <= 8'hC0; 15'h2047: d <= 8'hC0;
                15'h2048: d <= 8'hC0; 15'h2049: d <= 8'hC0; 15'h204A: d <= 8'hC0; 15'h204B: d <= 8'hC0;
                15'h204C: d <= 8'hC0; 15'h204D: d <= 8'hC0; 15'h204E: d <= 8'hC0; 15'h204F: d <= 8'hC0;
                15'h2050: d <= 8'hC0; 15'h2051: d <= 8'hC0; 15'h2052: d <= 8'hC0; 15'h2053: d <= 8'hC0;
                15'h2054: d <= 8'hC0; 15'h2055: d <= 8'hC0; 15'h2056: d <= 8'hC0; 15'h2057: d <= 8'hC0;
                15'h2058: d <= 8'hC0; 15'h2059: d <= 8'hC0; 15'h205A: d <= 8'hC0; 15'h205B: d <= 8'hC0;
                15'h205C: d <= 8'hC0; 15'h205D: d <= 8'hC0; 15'h205E: d <= 8'hC0; 15'h205F: d <= 8'hC0;
                15'h2060: d <= 8'hC0; 15'h2061: d <= 8'hC0; 15'h2062: d <= 8'hC0; 15'h2063: d <= 8'hC0;
                15'h2064: d <= 8'hC0; 15'h2065: d <= 8'hC0; 15'h2066: d <= 8'hC0; 15'h2067: d <= 8'hC0;
                15'h2068: d <= 8'hC0; 15'h2069: d <= 8'hC0; 15'h206A: d <= 8'hC0; 15'h206B: d <= 8'hC0;
                15'h206C: d <= 8'hC0; 15'h206D: d <= 8'hC0; 15'h206E: d <= 8'hC0; 15'h206F: d <= 8'hC0;
                15'h2070: d <= 8'hC0; 15'h2071: d <= 8'hC0; 15'h2072: d <= 8'hC0; 15'h2073: d <= 8'hC0;
                15'h2074: d <= 8'hC0; 15'h2075: d <= 8'hC0; 15'h2076: d <= 8'hC0; 15'h2077: d <= 8'hC0;
                15'h2078: d <= 8'hC0; 15'h2079: d <= 8'hC0; 15'h207A: d <= 8'hC0; 15'h207B: d <= 8'hC0;
                15'h207C: d <= 8'hC0; 15'h207D: d <= 8'hC0; 15'h207E: d <= 8'hC0; 15'h207F: d <= 8'hC0;
                15'h2080: d <= 8'hC0; 15'h2081: d <= 8'hC0; 15'h2082: d <= 8'hC0; 15'h2083: d <= 8'hC0;
                15'h2084: d <= 8'hC0; 15'h2085: d <= 8'hC0; 15'h2086: d <= 8'hC0; 15'h2087: d <= 8'hC0;
                15'h2088: d <= 8'hC0; 15'h2089: d <= 8'hC0; 15'h208A: d <= 8'hC0; 15'h208B: d <= 8'hC0;
                15'h208C: d <= 8'hC0; 15'h208D: d <= 8'hC0; 15'h208E: d <= 8'hC0; 15'h208F: d <= 8'hC0;
                15'h2090: d <= 8'hC0; 15'h2091: d <= 8'hC0; 15'h2092: d <= 8'hC0; 15'h2093: d <= 8'hC0;
                15'h2094: d <= 8'hC0; 15'h2095: d <= 8'hC0; 15'h2096: d <= 8'hC0; 15'h2097: d <= 8'hC0;
                15'h2098: d <= 8'hC0; 15'h2099: d <= 8'hC0; 15'h209A: d <= 8'hC0; 15'h209B: d <= 8'hC0;
                15'h209C: d <= 8'hC0; 15'h209D: d <= 8'hC0; 15'h209E: d <= 8'hC0; 15'h209F: d <= 8'hC0;
                15'h20A0: d <= 8'hC0; 15'h20A1: d <= 8'hC0; 15'h20A2: d <= 8'hC0; 15'h20A3: d <= 8'hC0;
                15'h20A4: d <= 8'hC0; 15'h20A5: d <= 8'hC0; 15'h20A6: d <= 8'hC0; 15'h20A7: d <= 8'hC0;
                15'h20A8: d <= 8'hC0; 15'h20A9: d <= 8'hC0; 15'h20AA: d <= 8'hC0; 15'h20AB: d <= 8'hC0;
                15'h20AC: d <= 8'hC0; 15'h20AD: d <= 8'hC0; 15'h20AE: d <= 8'hC0; 15'h20AF: d <= 8'hC0;
                15'h20B0: d <= 8'hC0; 15'h20B1: d <= 8'hC0; 15'h20B2: d <= 8'hC0; 15'h20B3: d <= 8'hC0;
                15'h20B4: d <= 8'hC0; 15'h20B5: d <= 8'hC0; 15'h20B6: d <= 8'hC0; 15'h20B7: d <= 8'hC0;
                15'h20B8: d <= 8'hC0; 15'h20B9: d <= 8'hC0; 15'h20BA: d <= 8'hC0; 15'h20BB: d <= 8'hC0;
                15'h20BC: d <= 8'hC0; 15'h20BD: d <= 8'hC0; 15'h20BE: d <= 8'hC0; 15'h20BF: d <= 8'hC0;
                15'h20C0: d <= 8'hC0; 15'h20C1: d <= 8'hC0; 15'h20C2: d <= 8'hC0; 15'h20C3: d <= 8'hC0;
                15'h20C4: d <= 8'hC0; 15'h20C5: d <= 8'hC0; 15'h20C6: d <= 8'hC0; 15'h20C7: d <= 8'hC0;
                15'h20C8: d <= 8'hC0; 15'h20C9: d <= 8'hC0; 15'h20CA: d <= 8'hC0; 15'h20CB: d <= 8'hC0;
                15'h20CC: d <= 8'hC0; 15'h20CD: d <= 8'hC0; 15'h20CE: d <= 8'hC0; 15'h20CF: d <= 8'hC0;
                15'h20D0: d <= 8'hC0; 15'h20D1: d <= 8'hC0; 15'h20D2: d <= 8'hC0; 15'h20D3: d <= 8'hC0;
                15'h20D4: d <= 8'hC0; 15'h20D5: d <= 8'hC0; 15'h20D6: d <= 8'hC0; 15'h20D7: d <= 8'hC0;
                15'h20D8: d <= 8'hC0; 15'h20D9: d <= 8'hC0; 15'h20DA: d <= 8'hC0; 15'h20DB: d <= 8'hC0;
                15'h20DC: d <= 8'hC0; 15'h20DD: d <= 8'hC0; 15'h20DE: d <= 8'hC0; 15'h20DF: d <= 8'hC0;
                15'h20E0: d <= 8'hC0; 15'h20E1: d <= 8'hC0; 15'h20E2: d <= 8'hC0; 15'h20E3: d <= 8'hC0;
                15'h20E4: d <= 8'hC0; 15'h20E5: d <= 8'hC0; 15'h20E6: d <= 8'hC0; 15'h20E7: d <= 8'hC0;
                15'h20E8: d <= 8'hC0; 15'h20E9: d <= 8'hC0; 15'h20EA: d <= 8'hC0; 15'h20EB: d <= 8'hC0;
                15'h20EC: d <= 8'hC0; 15'h20ED: d <= 8'hC0; 15'h20EE: d <= 8'hC0; 15'h20EF: d <= 8'hC0;
                15'h20F0: d <= 8'hC0; 15'h20F1: d <= 8'hC0; 15'h20F2: d <= 8'hC0; 15'h20F3: d <= 8'hC0;
                15'h20F4: d <= 8'hC0; 15'h20F5: d <= 8'hC0; 15'h20F6: d <= 8'hC0; 15'h20F7: d <= 8'hC0;
                15'h20F8: d <= 8'hC0; 15'h20F9: d <= 8'hC0; 15'h20FA: d <= 8'hC0; 15'h20FB: d <= 8'hC0;
                15'h20FC: d <= 8'hC0; 15'h20FD: d <= 8'hC0; 15'h20FE: d <= 8'hC0; 15'h20FF: d <= 8'hC0;
                15'h2100: d <= 8'hC0; 15'h2101: d <= 8'hC0; 15'h2102: d <= 8'hC0; 15'h2103: d <= 8'hC0;
                15'h2104: d <= 8'hC0; 15'h2105: d <= 8'hC0; 15'h2106: d <= 8'hC0; 15'h2107: d <= 8'hC0;
                15'h2108: d <= 8'hC0; 15'h2109: d <= 8'hC0; 15'h210A: d <= 8'hC0; 15'h210B: d <= 8'hC0;
                15'h210C: d <= 8'hC0; 15'h210D: d <= 8'hC0; 15'h210E: d <= 8'hC0; 15'h210F: d <= 8'hC0;
                15'h2110: d <= 8'hC0; 15'h2111: d <= 8'hC0; 15'h2112: d <= 8'hC0; 15'h2113: d <= 8'hC0;
                15'h2114: d <= 8'hC0; 15'h2115: d <= 8'hC0; 15'h2116: d <= 8'hC0; 15'h2117: d <= 8'hC0;
                15'h2118: d <= 8'hC0; 15'h2119: d <= 8'hC0; 15'h211A: d <= 8'hC0; 15'h211B: d <= 8'hC0;
                15'h211C: d <= 8'hC0; 15'h211D: d <= 8'hC0; 15'h211E: d <= 8'hC0; 15'h211F: d <= 8'hC0;
                15'h2120: d <= 8'hC0; 15'h2121: d <= 8'hC0; 15'h2122: d <= 8'hC0; 15'h2123: d <= 8'hC0;
                15'h2124: d <= 8'hC0; 15'h2125: d <= 8'hC0; 15'h2126: d <= 8'hC0; 15'h2127: d <= 8'hC0;
                15'h2128: d <= 8'hC0; 15'h2129: d <= 8'hC0; 15'h212A: d <= 8'hC0; 15'h212B: d <= 8'hC0;
                15'h212C: d <= 8'hC0; 15'h212D: d <= 8'hC0; 15'h212E: d <= 8'hC0; 15'h212F: d <= 8'hC0;
                15'h2130: d <= 8'hC0; 15'h2131: d <= 8'hC0; 15'h2132: d <= 8'hC0; 15'h2133: d <= 8'hC0;
                15'h2134: d <= 8'hC0; 15'h2135: d <= 8'hC0; 15'h2136: d <= 8'hC0; 15'h2137: d <= 8'hC0;
                15'h2138: d <= 8'hC0; 15'h2139: d <= 8'hC0; 15'h213A: d <= 8'hC0; 15'h213B: d <= 8'hC0;
                15'h213C: d <= 8'hC0; 15'h213D: d <= 8'hC0; 15'h213E: d <= 8'hC0; 15'h213F: d <= 8'hC0;
                15'h2140: d <= 8'hC0; 15'h2141: d <= 8'hC0; 15'h2142: d <= 8'hC0; 15'h2143: d <= 8'hC0;
                15'h2144: d <= 8'hC0; 15'h2145: d <= 8'hC0; 15'h2146: d <= 8'hC0; 15'h2147: d <= 8'hC0;
                15'h2148: d <= 8'hC0; 15'h2149: d <= 8'hC0; 15'h214A: d <= 8'hC0; 15'h214B: d <= 8'hC0;
                15'h214C: d <= 8'hC0; 15'h214D: d <= 8'hC0; 15'h214E: d <= 8'hC0; 15'h214F: d <= 8'hC0;
                15'h2150: d <= 8'hC0; 15'h2151: d <= 8'hC0; 15'h2152: d <= 8'hC0; 15'h2153: d <= 8'hC0;
                15'h2154: d <= 8'hC0; 15'h2155: d <= 8'hC0; 15'h2156: d <= 8'hC0; 15'h2157: d <= 8'hC0;
                15'h2158: d <= 8'hC0; 15'h2159: d <= 8'hC0; 15'h215A: d <= 8'hC0; 15'h215B: d <= 8'hC0;
                15'h215C: d <= 8'hC0; 15'h215D: d <= 8'hC0; 15'h215E: d <= 8'hC0; 15'h215F: d <= 8'hC0;
                15'h2160: d <= 8'hC0; 15'h2161: d <= 8'hC0; 15'h2162: d <= 8'hC0; 15'h2163: d <= 8'hC0;
                15'h2164: d <= 8'hC0; 15'h2165: d <= 8'hC0; 15'h2166: d <= 8'hC0; 15'h2167: d <= 8'hC0;
                15'h2168: d <= 8'hC0; 15'h2169: d <= 8'hC0; 15'h216A: d <= 8'hC0; 15'h216B: d <= 8'hC0;
                15'h216C: d <= 8'hC0; 15'h216D: d <= 8'hC0; 15'h216E: d <= 8'hC0; 15'h216F: d <= 8'hC0;
                15'h2170: d <= 8'hC0; 15'h2171: d <= 8'hC0; 15'h2172: d <= 8'hC0; 15'h2173: d <= 8'hC0;
                15'h2174: d <= 8'hC0; 15'h2175: d <= 8'hC0; 15'h2176: d <= 8'hC0; 15'h2177: d <= 8'hC0;
                15'h2178: d <= 8'hC0; 15'h2179: d <= 8'hC0; 15'h217A: d <= 8'hC0; 15'h217B: d <= 8'hC0;
                15'h217C: d <= 8'hC0; 15'h217D: d <= 8'hC0; 15'h217E: d <= 8'hC0; 15'h217F: d <= 8'hC0;
                15'h2180: d <= 8'hC0; 15'h2181: d <= 8'hC0; 15'h2182: d <= 8'hC0; 15'h2183: d <= 8'hC0;
                15'h2184: d <= 8'hC0; 15'h2185: d <= 8'hC0; 15'h2186: d <= 8'hC0; 15'h2187: d <= 8'hC0;
                15'h2188: d <= 8'hC0; 15'h2189: d <= 8'hC0; 15'h218A: d <= 8'hC0; 15'h218B: d <= 8'hC0;
                15'h218C: d <= 8'hC0; 15'h218D: d <= 8'hC0; 15'h218E: d <= 8'hC0; 15'h218F: d <= 8'hC0;
                15'h2190: d <= 8'hC0; 15'h2191: d <= 8'hC0; 15'h2192: d <= 8'hC0; 15'h2193: d <= 8'hC0;
                15'h2194: d <= 8'hC0; 15'h2195: d <= 8'hC0; 15'h2196: d <= 8'hC0; 15'h2197: d <= 8'hC0;
                15'h2198: d <= 8'hC0; 15'h2199: d <= 8'hC0; 15'h219A: d <= 8'hC0; 15'h219B: d <= 8'hC0;
                15'h219C: d <= 8'hC0; 15'h219D: d <= 8'hC0; 15'h219E: d <= 8'hC0; 15'h219F: d <= 8'hC0;
                15'h21A0: d <= 8'hC0; 15'h21A1: d <= 8'hC0; 15'h21A2: d <= 8'hC0; 15'h21A3: d <= 8'hC0;
                15'h21A4: d <= 8'hC0; 15'h21A5: d <= 8'hC0; 15'h21A6: d <= 8'hC0; 15'h21A7: d <= 8'hC0;
                15'h21A8: d <= 8'hC0; 15'h21A9: d <= 8'hC0; 15'h21AA: d <= 8'hC0; 15'h21AB: d <= 8'hC0;
                15'h21AC: d <= 8'hC0; 15'h21AD: d <= 8'hC0; 15'h21AE: d <= 8'hC0; 15'h21AF: d <= 8'hC0;
                15'h21B0: d <= 8'hC0; 15'h21B1: d <= 8'hC0; 15'h21B2: d <= 8'hC0; 15'h21B3: d <= 8'hC0;
                15'h21B4: d <= 8'hC0; 15'h21B5: d <= 8'hC0; 15'h21B6: d <= 8'hC0; 15'h21B7: d <= 8'hC0;
                15'h21B8: d <= 8'hC0; 15'h21B9: d <= 8'hC0; 15'h21BA: d <= 8'hC0; 15'h21BB: d <= 8'hC0;
                15'h21BC: d <= 8'hC0; 15'h21BD: d <= 8'hC0; 15'h21BE: d <= 8'hC0; 15'h21BF: d <= 8'hC0;
                15'h21C0: d <= 8'hC0; 15'h21C1: d <= 8'hC0; 15'h21C2: d <= 8'hC0; 15'h21C3: d <= 8'hC0;
                15'h21C4: d <= 8'hC0; 15'h21C5: d <= 8'hC0; 15'h21C6: d <= 8'hC0; 15'h21C7: d <= 8'hC0;
                15'h21C8: d <= 8'hC0; 15'h21C9: d <= 8'hC0; 15'h21CA: d <= 8'hC0; 15'h21CB: d <= 8'hC0;
                15'h21CC: d <= 8'hC0; 15'h21CD: d <= 8'hC0; 15'h21CE: d <= 8'hC0; 15'h21CF: d <= 8'hC0;
                15'h21D0: d <= 8'hC0; 15'h21D1: d <= 8'hC0; 15'h21D2: d <= 8'hC0; 15'h21D3: d <= 8'hC0;
                15'h21D4: d <= 8'hC0; 15'h21D5: d <= 8'hC0; 15'h21D6: d <= 8'hC0; 15'h21D7: d <= 8'hC0;
                15'h21D8: d <= 8'hC0; 15'h21D9: d <= 8'hC0; 15'h21DA: d <= 8'hC0; 15'h21DB: d <= 8'hC0;
                15'h21DC: d <= 8'hC0; 15'h21DD: d <= 8'hC0; 15'h21DE: d <= 8'hC0; 15'h21DF: d <= 8'hC0;
                15'h21E0: d <= 8'hC0; 15'h21E1: d <= 8'hC0; 15'h21E2: d <= 8'hC0; 15'h21E3: d <= 8'hC0;
                15'h21E4: d <= 8'hC0; 15'h21E5: d <= 8'hC0; 15'h21E6: d <= 8'hC0; 15'h21E7: d <= 8'hC0;
                15'h21E8: d <= 8'hC0; 15'h21E9: d <= 8'hC0; 15'h21EA: d <= 8'hC0; 15'h21EB: d <= 8'hC0;
                15'h21EC: d <= 8'hC0; 15'h21ED: d <= 8'hC0; 15'h21EE: d <= 8'hC0; 15'h21EF: d <= 8'hC0;
                15'h21F0: d <= 8'hC0; 15'h21F1: d <= 8'hC0; 15'h21F2: d <= 8'hC0; 15'h21F3: d <= 8'hC0;
                15'h21F4: d <= 8'hC0; 15'h21F5: d <= 8'hC0; 15'h21F6: d <= 8'hC0; 15'h21F7: d <= 8'hC0;
                15'h21F8: d <= 8'hC0; 15'h21F9: d <= 8'hC0; 15'h21FA: d <= 8'hC0; 15'h21FB: d <= 8'hC0;
                15'h21FC: d <= 8'hC0; 15'h21FD: d <= 8'hC0; 15'h21FE: d <= 8'hC0; 15'h21FF: d <= 8'hC0;
                15'h2200: d <= 8'hC0; 15'h2201: d <= 8'hC0; 15'h2202: d <= 8'hC0; 15'h2203: d <= 8'hC0;
                15'h2204: d <= 8'hC0; 15'h2205: d <= 8'hC0; 15'h2206: d <= 8'hC0; 15'h2207: d <= 8'hC0;
                15'h2208: d <= 8'hC0; 15'h2209: d <= 8'hC0; 15'h220A: d <= 8'hC0; 15'h220B: d <= 8'hC0;
                15'h220C: d <= 8'hC0; 15'h220D: d <= 8'hC0; 15'h220E: d <= 8'hC0; 15'h220F: d <= 8'hC0;
                15'h2210: d <= 8'hC0; 15'h2211: d <= 8'hC0; 15'h2212: d <= 8'hC0; 15'h2213: d <= 8'hC0;
                15'h2214: d <= 8'hC0; 15'h2215: d <= 8'hC0; 15'h2216: d <= 8'hC0; 15'h2217: d <= 8'hC0;
                15'h2218: d <= 8'hC0; 15'h2219: d <= 8'hC0; 15'h221A: d <= 8'hC0; 15'h221B: d <= 8'hC0;
                15'h221C: d <= 8'hC0; 15'h221D: d <= 8'hC0; 15'h221E: d <= 8'hC0; 15'h221F: d <= 8'hC0;
                15'h2220: d <= 8'hC0; 15'h2221: d <= 8'hC0; 15'h2222: d <= 8'hC0; 15'h2223: d <= 8'hC0;
                15'h2224: d <= 8'hC0; 15'h2225: d <= 8'hC0; 15'h2226: d <= 8'hC0; 15'h2227: d <= 8'hC0;
                15'h2228: d <= 8'hC0; 15'h2229: d <= 8'hC0; 15'h222A: d <= 8'hC0; 15'h222B: d <= 8'hC0;
                15'h222C: d <= 8'hC0; 15'h222D: d <= 8'hC0; 15'h222E: d <= 8'hC0; 15'h222F: d <= 8'hC0;
                15'h2230: d <= 8'hC0; 15'h2231: d <= 8'hC0; 15'h2232: d <= 8'hC0; 15'h2233: d <= 8'hC0;
                15'h2234: d <= 8'hC0; 15'h2235: d <= 8'hC0; 15'h2236: d <= 8'hC0; 15'h2237: d <= 8'hC0;
                15'h2238: d <= 8'hC0; 15'h2239: d <= 8'hC0; 15'h223A: d <= 8'hC0; 15'h223B: d <= 8'hC0;
                15'h223C: d <= 8'hC0; 15'h223D: d <= 8'hC0; 15'h223E: d <= 8'hC0; 15'h223F: d <= 8'hC0;
                15'h2240: d <= 8'hC0; 15'h2241: d <= 8'hC0; 15'h2242: d <= 8'hC0; 15'h2243: d <= 8'hC0;
                15'h2244: d <= 8'hC0; 15'h2245: d <= 8'hC0; 15'h2246: d <= 8'hC0; 15'h2247: d <= 8'hC0;
                15'h2248: d <= 8'hC0; 15'h2249: d <= 8'hC0; 15'h224A: d <= 8'hC0; 15'h224B: d <= 8'hC0;
                15'h224C: d <= 8'hC0; 15'h224D: d <= 8'hC0; 15'h224E: d <= 8'hC0; 15'h224F: d <= 8'hC0;
                15'h2250: d <= 8'hC0; 15'h2251: d <= 8'hC0; 15'h2252: d <= 8'hC0; 15'h2253: d <= 8'hC0;
                15'h2254: d <= 8'hC0; 15'h2255: d <= 8'hC0; 15'h2256: d <= 8'hC0; 15'h2257: d <= 8'hC0;
                15'h2258: d <= 8'hC0; 15'h2259: d <= 8'hC0; 15'h225A: d <= 8'hC0; 15'h225B: d <= 8'hC0;
                15'h225C: d <= 8'hC0; 15'h225D: d <= 8'hC0; 15'h225E: d <= 8'hC0; 15'h225F: d <= 8'hC0;
                15'h2260: d <= 8'hC0; 15'h2261: d <= 8'hC0; 15'h2262: d <= 8'hC0; 15'h2263: d <= 8'hC0;
                15'h2264: d <= 8'hC0; 15'h2265: d <= 8'hC0; 15'h2266: d <= 8'hC0; 15'h2267: d <= 8'hC0;
                15'h2268: d <= 8'hC0; 15'h2269: d <= 8'hC0; 15'h226A: d <= 8'hC0; 15'h226B: d <= 8'hC0;
                15'h226C: d <= 8'hC0; 15'h226D: d <= 8'hC0; 15'h226E: d <= 8'hC0; 15'h226F: d <= 8'hC0;
                15'h2270: d <= 8'hC0; 15'h2271: d <= 8'hC0; 15'h2272: d <= 8'hC0; 15'h2273: d <= 8'hC0;
                15'h2274: d <= 8'hC0; 15'h2275: d <= 8'hC0; 15'h2276: d <= 8'hC0; 15'h2277: d <= 8'hC0;
                15'h2278: d <= 8'hC0; 15'h2279: d <= 8'hC0; 15'h227A: d <= 8'hC0; 15'h227B: d <= 8'hC0;
                15'h227C: d <= 8'hC0; 15'h227D: d <= 8'hC0; 15'h227E: d <= 8'hC0; 15'h227F: d <= 8'hC0;
                15'h2280: d <= 8'hC0; 15'h2281: d <= 8'hC0; 15'h2282: d <= 8'hC0; 15'h2283: d <= 8'hC0;
                15'h2284: d <= 8'hC0; 15'h2285: d <= 8'hC0; 15'h2286: d <= 8'hC0; 15'h2287: d <= 8'hC0;
                15'h2288: d <= 8'hC0; 15'h2289: d <= 8'hC0; 15'h228A: d <= 8'hC0; 15'h228B: d <= 8'hC0;
                15'h228C: d <= 8'hC0; 15'h228D: d <= 8'hC0; 15'h228E: d <= 8'hC0; 15'h228F: d <= 8'hC0;
                15'h2290: d <= 8'hC0; 15'h2291: d <= 8'hC0; 15'h2292: d <= 8'hC0; 15'h2293: d <= 8'hC0;
                15'h2294: d <= 8'hC0; 15'h2295: d <= 8'hC0; 15'h2296: d <= 8'hC0; 15'h2297: d <= 8'hC0;
                15'h2298: d <= 8'hC0; 15'h2299: d <= 8'hC0; 15'h229A: d <= 8'hC0; 15'h229B: d <= 8'hC0;
                15'h229C: d <= 8'hC0; 15'h229D: d <= 8'hC0; 15'h229E: d <= 8'hC0; 15'h229F: d <= 8'hC0;
                15'h22A0: d <= 8'hC0; 15'h22A1: d <= 8'hC0; 15'h22A2: d <= 8'hC0; 15'h22A3: d <= 8'hC0;
                15'h22A4: d <= 8'hC0; 15'h22A5: d <= 8'hC0; 15'h22A6: d <= 8'hC0; 15'h22A7: d <= 8'hC0;
                15'h22A8: d <= 8'hC0; 15'h22A9: d <= 8'hC0; 15'h22AA: d <= 8'hC0; 15'h22AB: d <= 8'hC0;
                15'h22AC: d <= 8'hC0; 15'h22AD: d <= 8'hC0; 15'h22AE: d <= 8'hC0; 15'h22AF: d <= 8'hC0;
                15'h22B0: d <= 8'hC0; 15'h22B1: d <= 8'hC0; 15'h22B2: d <= 8'hC0; 15'h22B3: d <= 8'hC0;
                15'h22B4: d <= 8'hC0; 15'h22B5: d <= 8'hC0; 15'h22B6: d <= 8'hC0; 15'h22B7: d <= 8'hC0;
                15'h22B8: d <= 8'hC0; 15'h22B9: d <= 8'hC0; 15'h22BA: d <= 8'hC0; 15'h22BB: d <= 8'hC0;
                15'h22BC: d <= 8'hC0; 15'h22BD: d <= 8'hC0; 15'h22BE: d <= 8'hC0; 15'h22BF: d <= 8'hC0;
                15'h22C0: d <= 8'hC0; 15'h22C1: d <= 8'hC0; 15'h22C2: d <= 8'hC0; 15'h22C3: d <= 8'hC0;
                15'h22C4: d <= 8'hC0; 15'h22C5: d <= 8'hC0; 15'h22C6: d <= 8'hC0; 15'h22C7: d <= 8'hC0;
                15'h22C8: d <= 8'hC0; 15'h22C9: d <= 8'hC0; 15'h22CA: d <= 8'hC0; 15'h22CB: d <= 8'hC0;
                15'h22CC: d <= 8'hC0; 15'h22CD: d <= 8'hC0; 15'h22CE: d <= 8'hC0; 15'h22CF: d <= 8'hC0;
                15'h22D0: d <= 8'hC0; 15'h22D1: d <= 8'hC0; 15'h22D2: d <= 8'hC0; 15'h22D3: d <= 8'hC0;
                15'h22D4: d <= 8'hC0; 15'h22D5: d <= 8'hC0; 15'h22D6: d <= 8'hC0; 15'h22D7: d <= 8'hC0;
                15'h22D8: d <= 8'hC0; 15'h22D9: d <= 8'hC0; 15'h22DA: d <= 8'hC0; 15'h22DB: d <= 8'hC0;
                15'h22DC: d <= 8'hC0; 15'h22DD: d <= 8'hC0; 15'h22DE: d <= 8'hC0; 15'h22DF: d <= 8'hC0;
                15'h22E0: d <= 8'hC0; 15'h22E1: d <= 8'hC0; 15'h22E2: d <= 8'hC0; 15'h22E3: d <= 8'hC0;
                15'h22E4: d <= 8'hC0; 15'h22E5: d <= 8'hC0; 15'h22E6: d <= 8'hC0; 15'h22E7: d <= 8'hC0;
                15'h22E8: d <= 8'hC0; 15'h22E9: d <= 8'hC0; 15'h22EA: d <= 8'hC0; 15'h22EB: d <= 8'hC0;
                15'h22EC: d <= 8'hC0; 15'h22ED: d <= 8'hC0; 15'h22EE: d <= 8'hC0; 15'h22EF: d <= 8'hC0;
                15'h22F0: d <= 8'hC0; 15'h22F1: d <= 8'hC0; 15'h22F2: d <= 8'hC0; 15'h22F3: d <= 8'hC0;
                15'h22F4: d <= 8'hC0; 15'h22F5: d <= 8'hC0; 15'h22F6: d <= 8'hC0; 15'h22F7: d <= 8'hC0;
                15'h22F8: d <= 8'hC0; 15'h22F9: d <= 8'hC0; 15'h22FA: d <= 8'hC0; 15'h22FB: d <= 8'hC0;
                15'h22FC: d <= 8'hC0; 15'h22FD: d <= 8'hC0; 15'h22FE: d <= 8'hC0; 15'h22FF: d <= 8'hC0;
                15'h2300: d <= 8'hC0; 15'h2301: d <= 8'hC0; 15'h2302: d <= 8'hC0; 15'h2303: d <= 8'hC0;
                15'h2304: d <= 8'hC0; 15'h2305: d <= 8'hC0; 15'h2306: d <= 8'hC0; 15'h2307: d <= 8'hC0;
                15'h2308: d <= 8'hC0; 15'h2309: d <= 8'hC0; 15'h230A: d <= 8'hC0; 15'h230B: d <= 8'hC0;
                15'h230C: d <= 8'hC0; 15'h230D: d <= 8'hC0; 15'h230E: d <= 8'hC0; 15'h230F: d <= 8'hC0;
                15'h2310: d <= 8'hC0; 15'h2311: d <= 8'hC0; 15'h2312: d <= 8'hC0; 15'h2313: d <= 8'hC0;
                15'h2314: d <= 8'hC0; 15'h2315: d <= 8'hC0; 15'h2316: d <= 8'hC0; 15'h2317: d <= 8'hC0;
                15'h2318: d <= 8'hC0; 15'h2319: d <= 8'hC0; 15'h231A: d <= 8'hC0; 15'h231B: d <= 8'hC0;
                15'h231C: d <= 8'hC0; 15'h231D: d <= 8'hC0; 15'h231E: d <= 8'hC0; 15'h231F: d <= 8'hC0;
                15'h2320: d <= 8'hC0; 15'h2321: d <= 8'hC0; 15'h2322: d <= 8'hC0; 15'h2323: d <= 8'hC0;
                15'h2324: d <= 8'hC0; 15'h2325: d <= 8'hC0; 15'h2326: d <= 8'hC0; 15'h2327: d <= 8'hC0;
                15'h2328: d <= 8'hC0; 15'h2329: d <= 8'hC0; 15'h232A: d <= 8'hC0; 15'h232B: d <= 8'hC0;
                15'h232C: d <= 8'hC0; 15'h232D: d <= 8'hC0; 15'h232E: d <= 8'hC0; 15'h232F: d <= 8'hC0;
                15'h2330: d <= 8'hC0; 15'h2331: d <= 8'hC0; 15'h2332: d <= 8'hC0; 15'h2333: d <= 8'hC0;
                15'h2334: d <= 8'hC0; 15'h2335: d <= 8'hC0; 15'h2336: d <= 8'hC0; 15'h2337: d <= 8'hC0;
                15'h2338: d <= 8'hC0; 15'h2339: d <= 8'hC0; 15'h233A: d <= 8'hC0; 15'h233B: d <= 8'hC0;
                15'h233C: d <= 8'hC0; 15'h233D: d <= 8'hC0; 15'h233E: d <= 8'hC0; 15'h233F: d <= 8'hC0;
                15'h2340: d <= 8'hC0; 15'h2341: d <= 8'hC0; 15'h2342: d <= 8'hC0; 15'h2343: d <= 8'hC0;
                15'h2344: d <= 8'hC0; 15'h2345: d <= 8'hC0; 15'h2346: d <= 8'hC0; 15'h2347: d <= 8'hC0;
                15'h2348: d <= 8'hC0; 15'h2349: d <= 8'hC0; 15'h234A: d <= 8'hC0; 15'h234B: d <= 8'hC0;
                15'h234C: d <= 8'hC0; 15'h234D: d <= 8'hC0; 15'h234E: d <= 8'hC0; 15'h234F: d <= 8'hC0;
                15'h2350: d <= 8'hC0; 15'h2351: d <= 8'hC0; 15'h2352: d <= 8'hC0; 15'h2353: d <= 8'hC0;
                15'h2354: d <= 8'hC0; 15'h2355: d <= 8'hC0; 15'h2356: d <= 8'hC0; 15'h2357: d <= 8'hC0;
                15'h2358: d <= 8'hC0; 15'h2359: d <= 8'hC0; 15'h235A: d <= 8'hC0; 15'h235B: d <= 8'hC0;
                15'h235C: d <= 8'hC0; 15'h235D: d <= 8'hC0; 15'h235E: d <= 8'hC0; 15'h235F: d <= 8'hC0;
                15'h2360: d <= 8'hC0; 15'h2361: d <= 8'hC0; 15'h2362: d <= 8'hC0; 15'h2363: d <= 8'hC0;
                15'h2364: d <= 8'hC0; 15'h2365: d <= 8'hC0; 15'h2366: d <= 8'hC0; 15'h2367: d <= 8'hC0;
                15'h2368: d <= 8'hC0; 15'h2369: d <= 8'hC0; 15'h236A: d <= 8'hC0; 15'h236B: d <= 8'hC0;
                15'h236C: d <= 8'hC0; 15'h236D: d <= 8'hC0; 15'h236E: d <= 8'hC0; 15'h236F: d <= 8'hC0;
                15'h2370: d <= 8'hC0; 15'h2371: d <= 8'hC0; 15'h2372: d <= 8'hC0; 15'h2373: d <= 8'hC0;
                15'h2374: d <= 8'hC0; 15'h2375: d <= 8'hC0; 15'h2376: d <= 8'hC0; 15'h2377: d <= 8'hC0;
                15'h2378: d <= 8'hC0; 15'h2379: d <= 8'hC0; 15'h237A: d <= 8'hC0; 15'h237B: d <= 8'hC0;
                15'h237C: d <= 8'hC0; 15'h237D: d <= 8'hC0; 15'h237E: d <= 8'hC0; 15'h237F: d <= 8'hC0;
                15'h2380: d <= 8'hC0; 15'h2381: d <= 8'hC0; 15'h2382: d <= 8'hC0; 15'h2383: d <= 8'hC0;
                15'h2384: d <= 8'hC0; 15'h2385: d <= 8'hC0; 15'h2386: d <= 8'hC0; 15'h2387: d <= 8'hC0;
                15'h2388: d <= 8'hC0; 15'h2389: d <= 8'hC0; 15'h238A: d <= 8'hC0; 15'h238B: d <= 8'hC0;
                15'h238C: d <= 8'hC0; 15'h238D: d <= 8'hC0; 15'h238E: d <= 8'hC0; 15'h238F: d <= 8'hC0;
                15'h2390: d <= 8'hC0; 15'h2391: d <= 8'hC0; 15'h2392: d <= 8'hC0; 15'h2393: d <= 8'hC0;
                15'h2394: d <= 8'hC0; 15'h2395: d <= 8'hC0; 15'h2396: d <= 8'hC0; 15'h2397: d <= 8'hC0;
                15'h2398: d <= 8'hC0; 15'h2399: d <= 8'hC0; 15'h239A: d <= 8'hC0; 15'h239B: d <= 8'hC0;
                15'h239C: d <= 8'hC0; 15'h239D: d <= 8'hC0; 15'h239E: d <= 8'hC0; 15'h239F: d <= 8'hC0;
                15'h23A0: d <= 8'hC0; 15'h23A1: d <= 8'hC0; 15'h23A2: d <= 8'hC0; 15'h23A3: d <= 8'hC0;
                15'h23A4: d <= 8'hC0; 15'h23A5: d <= 8'hC0; 15'h23A6: d <= 8'hC0; 15'h23A7: d <= 8'hC0;
                15'h23A8: d <= 8'hC0; 15'h23A9: d <= 8'hC0; 15'h23AA: d <= 8'hC0; 15'h23AB: d <= 8'hC0;
                15'h23AC: d <= 8'hC0; 15'h23AD: d <= 8'hC0; 15'h23AE: d <= 8'hC0; 15'h23AF: d <= 8'hC0;
                15'h23B0: d <= 8'hC0; 15'h23B1: d <= 8'hC0; 15'h23B2: d <= 8'hC0; 15'h23B3: d <= 8'hC0;
                15'h23B4: d <= 8'hC0; 15'h23B5: d <= 8'hC0; 15'h23B6: d <= 8'hC0; 15'h23B7: d <= 8'hC0;
                15'h23B8: d <= 8'hC0; 15'h23B9: d <= 8'hC0; 15'h23BA: d <= 8'hC0; 15'h23BB: d <= 8'hC0;
                15'h23BC: d <= 8'hC0; 15'h23BD: d <= 8'hC0; 15'h23BE: d <= 8'hC0; 15'h23BF: d <= 8'hC0;
                15'h23C0: d <= 8'hC0; 15'h23C1: d <= 8'hC0; 15'h23C2: d <= 8'hC0; 15'h23C3: d <= 8'hC0;
                15'h23C4: d <= 8'hC0; 15'h23C5: d <= 8'hC0; 15'h23C6: d <= 8'hC0; 15'h23C7: d <= 8'hC0;
                15'h23C8: d <= 8'hC0; 15'h23C9: d <= 8'hC0; 15'h23CA: d <= 8'hC0; 15'h23CB: d <= 8'hC0;
                15'h23CC: d <= 8'hC0; 15'h23CD: d <= 8'hC0; 15'h23CE: d <= 8'hC0; 15'h23CF: d <= 8'hC0;
                15'h23D0: d <= 8'hC0; 15'h23D1: d <= 8'hC0; 15'h23D2: d <= 8'hC0; 15'h23D3: d <= 8'hC0;
                15'h23D4: d <= 8'hC0; 15'h23D5: d <= 8'hC0; 15'h23D6: d <= 8'hC0; 15'h23D7: d <= 8'hC0;
                15'h23D8: d <= 8'hC0; 15'h23D9: d <= 8'hC0; 15'h23DA: d <= 8'hC0; 15'h23DB: d <= 8'hC0;
                15'h23DC: d <= 8'hC0; 15'h23DD: d <= 8'hC0; 15'h23DE: d <= 8'hC0; 15'h23DF: d <= 8'hC0;
                15'h23E0: d <= 8'hC0; 15'h23E1: d <= 8'hC0; 15'h23E2: d <= 8'hC0; 15'h23E3: d <= 8'hC0;
                15'h23E4: d <= 8'hC0; 15'h23E5: d <= 8'hC0; 15'h23E6: d <= 8'hC0; 15'h23E7: d <= 8'hC0;
                15'h23E8: d <= 8'hC0; 15'h23E9: d <= 8'hC0; 15'h23EA: d <= 8'hC0; 15'h23EB: d <= 8'hC0;
                15'h23EC: d <= 8'hC0; 15'h23ED: d <= 8'hC0; 15'h23EE: d <= 8'hC0; 15'h23EF: d <= 8'hC0;
                15'h23F0: d <= 8'hC0; 15'h23F1: d <= 8'hC0; 15'h23F2: d <= 8'hC0; 15'h23F3: d <= 8'hC0;
                15'h23F4: d <= 8'hC0; 15'h23F5: d <= 8'hC0; 15'h23F6: d <= 8'hC0; 15'h23F7: d <= 8'hC0;
                15'h23F8: d <= 8'hC0; 15'h23F9: d <= 8'hC0; 15'h23FA: d <= 8'hC0; 15'h23FB: d <= 8'hC0;
                15'h23FC: d <= 8'hC0; 15'h23FD: d <= 8'hC0; 15'h23FE: d <= 8'hC0; 15'h23FF: d <= 8'hC0;
                15'h2400: d <= 8'hC0; 15'h2401: d <= 8'hC0; 15'h2402: d <= 8'hC0; 15'h2403: d <= 8'hC0;
                15'h2404: d <= 8'hC0; 15'h2405: d <= 8'hC0; 15'h2406: d <= 8'hC0; 15'h2407: d <= 8'hC0;
                15'h2408: d <= 8'hC0; 15'h2409: d <= 8'hC0; 15'h240A: d <= 8'hC0; 15'h240B: d <= 8'hC0;
                15'h240C: d <= 8'hC0; 15'h240D: d <= 8'hC0; 15'h240E: d <= 8'hC0; 15'h240F: d <= 8'hC0;
                15'h2410: d <= 8'hC0; 15'h2411: d <= 8'hC0; 15'h2412: d <= 8'hC0; 15'h2413: d <= 8'hC0;
                15'h2414: d <= 8'hC0; 15'h2415: d <= 8'hC0; 15'h2416: d <= 8'hC0; 15'h2417: d <= 8'hC0;
                15'h2418: d <= 8'hC0; 15'h2419: d <= 8'hC0; 15'h241A: d <= 8'hC0; 15'h241B: d <= 8'hC0;
                15'h241C: d <= 8'hC0; 15'h241D: d <= 8'hC0; 15'h241E: d <= 8'hC0; 15'h241F: d <= 8'hC0;
                15'h2420: d <= 8'hC0; 15'h2421: d <= 8'hC0; 15'h2422: d <= 8'hC0; 15'h2423: d <= 8'hC0;
                15'h2424: d <= 8'hC0; 15'h2425: d <= 8'hC0; 15'h2426: d <= 8'hC0; 15'h2427: d <= 8'hC0;
                15'h2428: d <= 8'hC0; 15'h2429: d <= 8'hC0; 15'h242A: d <= 8'hC0; 15'h242B: d <= 8'hC0;
                15'h242C: d <= 8'hC0; 15'h242D: d <= 8'hC0; 15'h242E: d <= 8'hC0; 15'h242F: d <= 8'hC0;
                15'h2430: d <= 8'hC0; 15'h2431: d <= 8'hC0; 15'h2432: d <= 8'hC0; 15'h2433: d <= 8'hC0;
                15'h2434: d <= 8'hC0; 15'h2435: d <= 8'hC0; 15'h2436: d <= 8'hC0; 15'h2437: d <= 8'hC0;
                15'h2438: d <= 8'hC0; 15'h2439: d <= 8'hC0; 15'h243A: d <= 8'hC0; 15'h243B: d <= 8'hC0;
                15'h243C: d <= 8'hC0; 15'h243D: d <= 8'hC0; 15'h243E: d <= 8'hC0; 15'h243F: d <= 8'hC0;
                15'h2440: d <= 8'hC0; 15'h2441: d <= 8'hC0; 15'h2442: d <= 8'hC0; 15'h2443: d <= 8'hC0;
                15'h2444: d <= 8'hC0; 15'h2445: d <= 8'hC0; 15'h2446: d <= 8'hC0; 15'h2447: d <= 8'hC0;
                15'h2448: d <= 8'hC0; 15'h2449: d <= 8'hC0; 15'h244A: d <= 8'hC0; 15'h244B: d <= 8'hC0;
                15'h244C: d <= 8'hC0; 15'h244D: d <= 8'hC0; 15'h244E: d <= 8'hC0; 15'h244F: d <= 8'hC0;
                15'h2450: d <= 8'hC0; 15'h2451: d <= 8'hC0; 15'h2452: d <= 8'hC0; 15'h2453: d <= 8'hC0;
                15'h2454: d <= 8'hC0; 15'h2455: d <= 8'hC0; 15'h2456: d <= 8'hC0; 15'h2457: d <= 8'hC0;
                15'h2458: d <= 8'hC0; 15'h2459: d <= 8'hC0; 15'h245A: d <= 8'hC0; 15'h245B: d <= 8'hC0;
                15'h245C: d <= 8'hC0; 15'h245D: d <= 8'hC0; 15'h245E: d <= 8'hC0; 15'h245F: d <= 8'hC0;
                15'h2460: d <= 8'hC0; 15'h2461: d <= 8'hC0; 15'h2462: d <= 8'hC0; 15'h2463: d <= 8'hC0;
                15'h2464: d <= 8'hC0; 15'h2465: d <= 8'hC0; 15'h2466: d <= 8'hC0; 15'h2467: d <= 8'hC0;
                15'h2468: d <= 8'hC0; 15'h2469: d <= 8'hC0; 15'h246A: d <= 8'hC0; 15'h246B: d <= 8'hC0;
                15'h246C: d <= 8'hC0; 15'h246D: d <= 8'hC0; 15'h246E: d <= 8'hC0; 15'h246F: d <= 8'hC0;
                15'h2470: d <= 8'hC0; 15'h2471: d <= 8'hC0; 15'h2472: d <= 8'hC0; 15'h2473: d <= 8'hC0;
                15'h2474: d <= 8'hC0; 15'h2475: d <= 8'hC0; 15'h2476: d <= 8'hC0; 15'h2477: d <= 8'hC0;
                15'h2478: d <= 8'hC0; 15'h2479: d <= 8'hC0; 15'h247A: d <= 8'hC0; 15'h247B: d <= 8'hC0;
                15'h247C: d <= 8'hC0; 15'h247D: d <= 8'hC0; 15'h247E: d <= 8'hC0; 15'h247F: d <= 8'hC0;
                15'h2480: d <= 8'hC0; 15'h2481: d <= 8'hC0; 15'h2482: d <= 8'hC0; 15'h2483: d <= 8'hC0;
                15'h2484: d <= 8'hC0; 15'h2485: d <= 8'hC0; 15'h2486: d <= 8'hC0; 15'h2487: d <= 8'hC0;
                15'h2488: d <= 8'hC0; 15'h2489: d <= 8'hC0; 15'h248A: d <= 8'hC0; 15'h248B: d <= 8'hC0;
                15'h248C: d <= 8'hC0; 15'h248D: d <= 8'hC0; 15'h248E: d <= 8'hC0; 15'h248F: d <= 8'hC0;
                15'h2490: d <= 8'hC0; 15'h2491: d <= 8'hC0; 15'h2492: d <= 8'hC0; 15'h2493: d <= 8'hC0;
                15'h2494: d <= 8'hC0; 15'h2495: d <= 8'hC0; 15'h2496: d <= 8'hC0; 15'h2497: d <= 8'hC0;
                15'h2498: d <= 8'hC0; 15'h2499: d <= 8'hC0; 15'h249A: d <= 8'hC0; 15'h249B: d <= 8'hC0;
                15'h249C: d <= 8'hC0; 15'h249D: d <= 8'hC0; 15'h249E: d <= 8'hC0; 15'h249F: d <= 8'hC0;
                15'h24A0: d <= 8'hC0; 15'h24A1: d <= 8'hC0; 15'h24A2: d <= 8'hC0; 15'h24A3: d <= 8'hC0;
                15'h24A4: d <= 8'hC0; 15'h24A5: d <= 8'hC0; 15'h24A6: d <= 8'hC0; 15'h24A7: d <= 8'hC0;
                15'h24A8: d <= 8'hC0; 15'h24A9: d <= 8'hC0; 15'h24AA: d <= 8'hC0; 15'h24AB: d <= 8'hC0;
                15'h24AC: d <= 8'hC0; 15'h24AD: d <= 8'hC0; 15'h24AE: d <= 8'hC0; 15'h24AF: d <= 8'hC0;
                15'h24B0: d <= 8'hC0; 15'h24B1: d <= 8'hC0; 15'h24B2: d <= 8'hC0; 15'h24B3: d <= 8'hC0;
                15'h24B4: d <= 8'hC0; 15'h24B5: d <= 8'hC0; 15'h24B6: d <= 8'hC0; 15'h24B7: d <= 8'hC0;
                15'h24B8: d <= 8'hC0; 15'h24B9: d <= 8'hC0; 15'h24BA: d <= 8'hC0; 15'h24BB: d <= 8'hC0;
                15'h24BC: d <= 8'hC0; 15'h24BD: d <= 8'hC0; 15'h24BE: d <= 8'hC0; 15'h24BF: d <= 8'hC0;
                15'h24C0: d <= 8'hC0; 15'h24C1: d <= 8'hC0; 15'h24C2: d <= 8'hC0; 15'h24C3: d <= 8'hC0;
                15'h24C4: d <= 8'hC0; 15'h24C5: d <= 8'hC0; 15'h24C6: d <= 8'hC0; 15'h24C7: d <= 8'hC0;
                15'h24C8: d <= 8'hC0; 15'h24C9: d <= 8'hC0; 15'h24CA: d <= 8'hC0; 15'h24CB: d <= 8'hC0;
                15'h24CC: d <= 8'hC0; 15'h24CD: d <= 8'hC0; 15'h24CE: d <= 8'hC0; 15'h24CF: d <= 8'hC0;
                15'h24D0: d <= 8'hC0; 15'h24D1: d <= 8'hC0; 15'h24D2: d <= 8'hC0; 15'h24D3: d <= 8'hC0;
                15'h24D4: d <= 8'hC0; 15'h24D5: d <= 8'hC0; 15'h24D6: d <= 8'hC0; 15'h24D7: d <= 8'hC0;
                15'h24D8: d <= 8'hC0; 15'h24D9: d <= 8'hC0; 15'h24DA: d <= 8'hC0; 15'h24DB: d <= 8'hC0;
                15'h24DC: d <= 8'hC0; 15'h24DD: d <= 8'hC0; 15'h24DE: d <= 8'hC0; 15'h24DF: d <= 8'hC0;
                15'h24E0: d <= 8'hC0; 15'h24E1: d <= 8'hC0; 15'h24E2: d <= 8'hC0; 15'h24E3: d <= 8'hC0;
                15'h24E4: d <= 8'hC0; 15'h24E5: d <= 8'hC0; 15'h24E6: d <= 8'hC0; 15'h24E7: d <= 8'hC0;
                15'h24E8: d <= 8'hC0; 15'h24E9: d <= 8'hC0; 15'h24EA: d <= 8'hC0; 15'h24EB: d <= 8'hC0;
                15'h24EC: d <= 8'hC0; 15'h24ED: d <= 8'hC0; 15'h24EE: d <= 8'hC0; 15'h24EF: d <= 8'hC0;
                15'h24F0: d <= 8'hC0; 15'h24F1: d <= 8'hC0; 15'h24F2: d <= 8'hC0; 15'h24F3: d <= 8'hC0;
                15'h24F4: d <= 8'hC0; 15'h24F5: d <= 8'hC0; 15'h24F6: d <= 8'hC0; 15'h24F7: d <= 8'hC0;
                15'h24F8: d <= 8'hC0; 15'h24F9: d <= 8'hC0; 15'h24FA: d <= 8'hC0; 15'h24FB: d <= 8'hC0;
                15'h24FC: d <= 8'hC0; 15'h24FD: d <= 8'hC0; 15'h24FE: d <= 8'hC0; 15'h24FF: d <= 8'hC0;
                15'h2500: d <= 8'hC0; 15'h2501: d <= 8'hC0; 15'h2502: d <= 8'hC0; 15'h2503: d <= 8'hC0;
                15'h2504: d <= 8'hC0; 15'h2505: d <= 8'hC0; 15'h2506: d <= 8'hC0; 15'h2507: d <= 8'hC0;
                15'h2508: d <= 8'hC0; 15'h2509: d <= 8'hC0; 15'h250A: d <= 8'hC0; 15'h250B: d <= 8'hC0;
                15'h250C: d <= 8'hC0; 15'h250D: d <= 8'hC0; 15'h250E: d <= 8'hC0; 15'h250F: d <= 8'hC0;
                15'h2510: d <= 8'hC0; 15'h2511: d <= 8'hC0; 15'h2512: d <= 8'hC0; 15'h2513: d <= 8'hC0;
                15'h2514: d <= 8'hC0; 15'h2515: d <= 8'hC0; 15'h2516: d <= 8'hC0; 15'h2517: d <= 8'hC0;
                15'h2518: d <= 8'hC0; 15'h2519: d <= 8'hC0; 15'h251A: d <= 8'hC0; 15'h251B: d <= 8'hC0;
                15'h251C: d <= 8'hC0; 15'h251D: d <= 8'hC0; 15'h251E: d <= 8'hC0; 15'h251F: d <= 8'hC0;
                15'h2520: d <= 8'hC0; 15'h2521: d <= 8'hC0; 15'h2522: d <= 8'hC0; 15'h2523: d <= 8'hC0;
                15'h2524: d <= 8'hC0; 15'h2525: d <= 8'hC0; 15'h2526: d <= 8'hC0; 15'h2527: d <= 8'hC0;
                15'h2528: d <= 8'hC0; 15'h2529: d <= 8'hC0; 15'h252A: d <= 8'hC0; 15'h252B: d <= 8'hC0;
                15'h252C: d <= 8'hC0; 15'h252D: d <= 8'hC0; 15'h252E: d <= 8'hC0; 15'h252F: d <= 8'hC0;
                15'h2530: d <= 8'hC0; 15'h2531: d <= 8'hC0; 15'h2532: d <= 8'hC0; 15'h2533: d <= 8'hC0;
                15'h2534: d <= 8'hC0; 15'h2535: d <= 8'hC0; 15'h2536: d <= 8'hC0; 15'h2537: d <= 8'hC0;
                15'h2538: d <= 8'hC0; 15'h2539: d <= 8'hC0; 15'h253A: d <= 8'hC0; 15'h253B: d <= 8'hC0;
                15'h253C: d <= 8'hC0; 15'h253D: d <= 8'hC0; 15'h253E: d <= 8'hC0; 15'h253F: d <= 8'hC0;
                15'h2540: d <= 8'hC0; 15'h2541: d <= 8'hC0; 15'h2542: d <= 8'hC0; 15'h2543: d <= 8'hC0;
                15'h2544: d <= 8'hC0; 15'h2545: d <= 8'hC0; 15'h2546: d <= 8'hC0; 15'h2547: d <= 8'hC0;
                15'h2548: d <= 8'hC0; 15'h2549: d <= 8'hC0; 15'h254A: d <= 8'hC0; 15'h254B: d <= 8'hC0;
                15'h254C: d <= 8'hC0; 15'h254D: d <= 8'hC0; 15'h254E: d <= 8'hC0; 15'h254F: d <= 8'hC0;
                15'h2550: d <= 8'hC0; 15'h2551: d <= 8'hC0; 15'h2552: d <= 8'hC0; 15'h2553: d <= 8'hC0;
                15'h2554: d <= 8'hC0; 15'h2555: d <= 8'hC0; 15'h2556: d <= 8'hC0; 15'h2557: d <= 8'hC0;
                15'h2558: d <= 8'hC0; 15'h2559: d <= 8'hC0; 15'h255A: d <= 8'hC0; 15'h255B: d <= 8'hC0;
                15'h255C: d <= 8'hC0; 15'h255D: d <= 8'hC0; 15'h255E: d <= 8'hC0; 15'h255F: d <= 8'hC0;
                15'h2560: d <= 8'hC0; 15'h2561: d <= 8'hC0; 15'h2562: d <= 8'hC0; 15'h2563: d <= 8'hC0;
                15'h2564: d <= 8'hC0; 15'h2565: d <= 8'hC0; 15'h2566: d <= 8'hC0; 15'h2567: d <= 8'hC0;
                15'h2568: d <= 8'hC0; 15'h2569: d <= 8'hC0; 15'h256A: d <= 8'hC0; 15'h256B: d <= 8'hC0;
                15'h256C: d <= 8'hC0; 15'h256D: d <= 8'hC0; 15'h256E: d <= 8'hC0; 15'h256F: d <= 8'hC0;
                15'h2570: d <= 8'hC0; 15'h2571: d <= 8'hC0; 15'h2572: d <= 8'hC0; 15'h2573: d <= 8'hC0;
                15'h2574: d <= 8'hC0; 15'h2575: d <= 8'hC0; 15'h2576: d <= 8'hC0; 15'h2577: d <= 8'hC0;
                15'h2578: d <= 8'hC0; 15'h2579: d <= 8'hC0; 15'h257A: d <= 8'hC0; 15'h257B: d <= 8'hC0;
                15'h257C: d <= 8'hC0; 15'h257D: d <= 8'hC0; 15'h257E: d <= 8'hC0; 15'h257F: d <= 8'hC0;
                15'h2580: d <= 8'hC0; 15'h2581: d <= 8'hC0; 15'h2582: d <= 8'hC0; 15'h2583: d <= 8'hC0;
                15'h2584: d <= 8'hC0; 15'h2585: d <= 8'hC0; 15'h2586: d <= 8'hC0; 15'h2587: d <= 8'hC0;
                15'h2588: d <= 8'hC0; 15'h2589: d <= 8'hC0; 15'h258A: d <= 8'hC0; 15'h258B: d <= 8'hC0;
                15'h258C: d <= 8'hC0; 15'h258D: d <= 8'hC0; 15'h258E: d <= 8'hC0; 15'h258F: d <= 8'hC0;
                15'h2590: d <= 8'hC0; 15'h2591: d <= 8'hC0; 15'h2592: d <= 8'hC0; 15'h2593: d <= 8'hC0;
                15'h2594: d <= 8'hC0; 15'h2595: d <= 8'hC0; 15'h2596: d <= 8'hC0; 15'h2597: d <= 8'hC0;
                15'h2598: d <= 8'hC0; 15'h2599: d <= 8'hC0; 15'h259A: d <= 8'hC0; 15'h259B: d <= 8'hC0;
                15'h259C: d <= 8'hC0; 15'h259D: d <= 8'hC0; 15'h259E: d <= 8'hC0; 15'h259F: d <= 8'hC0;
                15'h25A0: d <= 8'hC0; 15'h25A1: d <= 8'hC0; 15'h25A2: d <= 8'hC0; 15'h25A3: d <= 8'hC0;
                15'h25A4: d <= 8'hC0; 15'h25A5: d <= 8'hC0; 15'h25A6: d <= 8'hC0; 15'h25A7: d <= 8'hC0;
                15'h25A8: d <= 8'hC0; 15'h25A9: d <= 8'hC0; 15'h25AA: d <= 8'hC0; 15'h25AB: d <= 8'hC0;
                15'h25AC: d <= 8'hC0; 15'h25AD: d <= 8'hC0; 15'h25AE: d <= 8'hC0; 15'h25AF: d <= 8'hC0;
                15'h25B0: d <= 8'hC0; 15'h25B1: d <= 8'hC0; 15'h25B2: d <= 8'hC0; 15'h25B3: d <= 8'hC0;
                15'h25B4: d <= 8'hC0; 15'h25B5: d <= 8'hC0; 15'h25B6: d <= 8'hC0; 15'h25B7: d <= 8'hC0;
                15'h25B8: d <= 8'hC0; 15'h25B9: d <= 8'hC0; 15'h25BA: d <= 8'hC0; 15'h25BB: d <= 8'hC0;
                15'h25BC: d <= 8'hC0; 15'h25BD: d <= 8'hC0; 15'h25BE: d <= 8'hC0; 15'h25BF: d <= 8'hC0;
                15'h25C0: d <= 8'hC0; 15'h25C1: d <= 8'hC0; 15'h25C2: d <= 8'hC0; 15'h25C3: d <= 8'hC0;
                15'h25C4: d <= 8'hC0; 15'h25C5: d <= 8'hC0; 15'h25C6: d <= 8'hC0; 15'h25C7: d <= 8'hC0;
                15'h25C8: d <= 8'hC0; 15'h25C9: d <= 8'hC0; 15'h25CA: d <= 8'hC0; 15'h25CB: d <= 8'hC0;
                15'h25CC: d <= 8'hC0; 15'h25CD: d <= 8'hC0; 15'h25CE: d <= 8'hC0; 15'h25CF: d <= 8'hC0;
                15'h25D0: d <= 8'hC0; 15'h25D1: d <= 8'hC0; 15'h25D2: d <= 8'hC0; 15'h25D3: d <= 8'hC0;
                15'h25D4: d <= 8'hC0; 15'h25D5: d <= 8'hC0; 15'h25D6: d <= 8'hC0; 15'h25D7: d <= 8'hC0;
                15'h25D8: d <= 8'hC0; 15'h25D9: d <= 8'hC0; 15'h25DA: d <= 8'hC0; 15'h25DB: d <= 8'hC0;
                15'h25DC: d <= 8'hC0; 15'h25DD: d <= 8'hC0; 15'h25DE: d <= 8'hC0; 15'h25DF: d <= 8'hC0;
                15'h25E0: d <= 8'hC0; 15'h25E1: d <= 8'hC0; 15'h25E2: d <= 8'hC0; 15'h25E3: d <= 8'hC0;
                15'h25E4: d <= 8'hC0; 15'h25E5: d <= 8'hC0; 15'h25E6: d <= 8'hC0; 15'h25E7: d <= 8'hC0;
                15'h25E8: d <= 8'hC0; 15'h25E9: d <= 8'hC0; 15'h25EA: d <= 8'hC0; 15'h25EB: d <= 8'hC0;
                15'h25EC: d <= 8'hC0; 15'h25ED: d <= 8'hC0; 15'h25EE: d <= 8'hC0; 15'h25EF: d <= 8'hC0;
                15'h25F0: d <= 8'hC0; 15'h25F1: d <= 8'hC0; 15'h25F2: d <= 8'hC0; 15'h25F3: d <= 8'hC0;
                15'h25F4: d <= 8'hC0; 15'h25F5: d <= 8'hC0; 15'h25F6: d <= 8'hC0; 15'h25F7: d <= 8'hC0;
                15'h25F8: d <= 8'hC0; 15'h25F9: d <= 8'hC0; 15'h25FA: d <= 8'hC0; 15'h25FB: d <= 8'hC0;
                15'h25FC: d <= 8'hC0; 15'h25FD: d <= 8'hC0; 15'h25FE: d <= 8'hC0; 15'h25FF: d <= 8'hC0;
                15'h2600: d <= 8'hC0; 15'h2601: d <= 8'hC0; 15'h2602: d <= 8'hC0; 15'h2603: d <= 8'hC0;
                15'h2604: d <= 8'hC0; 15'h2605: d <= 8'hC0; 15'h2606: d <= 8'hC0; 15'h2607: d <= 8'hC0;
                15'h2608: d <= 8'hC0; 15'h2609: d <= 8'hC0; 15'h260A: d <= 8'hC0; 15'h260B: d <= 8'hC0;
                15'h260C: d <= 8'hC0; 15'h260D: d <= 8'hC0; 15'h260E: d <= 8'hC0; 15'h260F: d <= 8'hC0;
                15'h2610: d <= 8'hC0; 15'h2611: d <= 8'hC0; 15'h2612: d <= 8'hC0; 15'h2613: d <= 8'hC0;
                15'h2614: d <= 8'hC0; 15'h2615: d <= 8'hC0; 15'h2616: d <= 8'hC0; 15'h2617: d <= 8'hC0;
                15'h2618: d <= 8'hC0; 15'h2619: d <= 8'hC0; 15'h261A: d <= 8'hC0; 15'h261B: d <= 8'hC0;
                15'h261C: d <= 8'hC0; 15'h261D: d <= 8'hC0; 15'h261E: d <= 8'hC0; 15'h261F: d <= 8'hC0;
                15'h2620: d <= 8'hC0; 15'h2621: d <= 8'hC0; 15'h2622: d <= 8'hC0; 15'h2623: d <= 8'hC0;
                15'h2624: d <= 8'hC0; 15'h2625: d <= 8'hC0; 15'h2626: d <= 8'hC0; 15'h2627: d <= 8'hC0;
                15'h2628: d <= 8'hC0; 15'h2629: d <= 8'hC0; 15'h262A: d <= 8'hC0; 15'h262B: d <= 8'hC0;
                15'h262C: d <= 8'hC0; 15'h262D: d <= 8'hC0; 15'h262E: d <= 8'hC0; 15'h262F: d <= 8'hC0;
                15'h2630: d <= 8'hC0; 15'h2631: d <= 8'hC0; 15'h2632: d <= 8'hC0; 15'h2633: d <= 8'hC0;
                15'h2634: d <= 8'hC0; 15'h2635: d <= 8'hC0; 15'h2636: d <= 8'hC0; 15'h2637: d <= 8'hC0;
                15'h2638: d <= 8'hC0; 15'h2639: d <= 8'hC0; 15'h263A: d <= 8'hC0; 15'h263B: d <= 8'hC0;
                15'h263C: d <= 8'hC0; 15'h263D: d <= 8'hC0; 15'h263E: d <= 8'hC0; 15'h263F: d <= 8'hC0;
                15'h2640: d <= 8'hC0; 15'h2641: d <= 8'hC0; 15'h2642: d <= 8'hC0; 15'h2643: d <= 8'hC0;
                15'h2644: d <= 8'hC0; 15'h2645: d <= 8'hC0; 15'h2646: d <= 8'hC0; 15'h2647: d <= 8'hC0;
                15'h2648: d <= 8'hC0; 15'h2649: d <= 8'hC0; 15'h264A: d <= 8'hC0; 15'h264B: d <= 8'hC0;
                15'h264C: d <= 8'hC0; 15'h264D: d <= 8'hC0; 15'h264E: d <= 8'hC0; 15'h264F: d <= 8'hC0;
                15'h2650: d <= 8'hC0; 15'h2651: d <= 8'hC0; 15'h2652: d <= 8'hC0; 15'h2653: d <= 8'hC0;
                15'h2654: d <= 8'hC0; 15'h2655: d <= 8'hC0; 15'h2656: d <= 8'hC0; 15'h2657: d <= 8'hC0;
                15'h2658: d <= 8'hC0; 15'h2659: d <= 8'hC0; 15'h265A: d <= 8'hC0; 15'h265B: d <= 8'hC0;
                15'h265C: d <= 8'hC0; 15'h265D: d <= 8'hC0; 15'h265E: d <= 8'hC0; 15'h265F: d <= 8'hC0;
                15'h2660: d <= 8'hC0; 15'h2661: d <= 8'hC0; 15'h2662: d <= 8'hC0; 15'h2663: d <= 8'hC0;
                15'h2664: d <= 8'hC0; 15'h2665: d <= 8'hC0; 15'h2666: d <= 8'hC0; 15'h2667: d <= 8'hC0;
                15'h2668: d <= 8'hC0; 15'h2669: d <= 8'hC0; 15'h266A: d <= 8'hC0; 15'h266B: d <= 8'hC0;
                15'h266C: d <= 8'hC0; 15'h266D: d <= 8'hC0; 15'h266E: d <= 8'hC0; 15'h266F: d <= 8'hC0;
                15'h2670: d <= 8'hC0; 15'h2671: d <= 8'hC0; 15'h2672: d <= 8'hC0; 15'h2673: d <= 8'hC0;
                15'h2674: d <= 8'hC0; 15'h2675: d <= 8'hC0; 15'h2676: d <= 8'hC0; 15'h2677: d <= 8'hC0;
                15'h2678: d <= 8'hC0; 15'h2679: d <= 8'hC0; 15'h267A: d <= 8'hC0; 15'h267B: d <= 8'hC0;
                15'h267C: d <= 8'hC0; 15'h267D: d <= 8'hC0; 15'h267E: d <= 8'hC0; 15'h267F: d <= 8'hC0;
                15'h2680: d <= 8'hC0; 15'h2681: d <= 8'hC0; 15'h2682: d <= 8'hC0; 15'h2683: d <= 8'hC0;
                15'h2684: d <= 8'hC0; 15'h2685: d <= 8'hC0; 15'h2686: d <= 8'hC0; 15'h2687: d <= 8'hC0;
                15'h2688: d <= 8'hC0; 15'h2689: d <= 8'hC0; 15'h268A: d <= 8'hC0; 15'h268B: d <= 8'hC0;
                15'h268C: d <= 8'hC0; 15'h268D: d <= 8'hC0; 15'h268E: d <= 8'hC0; 15'h268F: d <= 8'hC0;
                15'h2690: d <= 8'hC0; 15'h2691: d <= 8'hC0; 15'h2692: d <= 8'hC0; 15'h2693: d <= 8'hC0;
                15'h2694: d <= 8'hC0; 15'h2695: d <= 8'hC0; 15'h2696: d <= 8'hC0; 15'h2697: d <= 8'hC0;
                15'h2698: d <= 8'hC0; 15'h2699: d <= 8'hC0; 15'h269A: d <= 8'hC0; 15'h269B: d <= 8'hC0;
                15'h269C: d <= 8'hC0; 15'h269D: d <= 8'hC0; 15'h269E: d <= 8'hC0; 15'h269F: d <= 8'hC0;
                15'h26A0: d <= 8'hC0; 15'h26A1: d <= 8'hC0; 15'h26A2: d <= 8'hC0; 15'h26A3: d <= 8'hC0;
                15'h26A4: d <= 8'hC0; 15'h26A5: d <= 8'hC0; 15'h26A6: d <= 8'hC0; 15'h26A7: d <= 8'hC0;
                15'h26A8: d <= 8'hC0; 15'h26A9: d <= 8'hC0; 15'h26AA: d <= 8'hC0; 15'h26AB: d <= 8'hC0;
                15'h26AC: d <= 8'hC0; 15'h26AD: d <= 8'hC0; 15'h26AE: d <= 8'hC0; 15'h26AF: d <= 8'hC0;
                15'h26B0: d <= 8'hC0; 15'h26B1: d <= 8'hC0; 15'h26B2: d <= 8'hC0; 15'h26B3: d <= 8'hC0;
                15'h26B4: d <= 8'hC0; 15'h26B5: d <= 8'hC0; 15'h26B6: d <= 8'hC0; 15'h26B7: d <= 8'hC0;
                15'h26B8: d <= 8'hC0; 15'h26B9: d <= 8'hC0; 15'h26BA: d <= 8'hC0; 15'h26BB: d <= 8'hC0;
                15'h26BC: d <= 8'hC0; 15'h26BD: d <= 8'hC0; 15'h26BE: d <= 8'hC0; 15'h26BF: d <= 8'hC0;
                15'h26C0: d <= 8'hC0; 15'h26C1: d <= 8'hC0; 15'h26C2: d <= 8'hC0; 15'h26C3: d <= 8'hC0;
                15'h26C4: d <= 8'hC0; 15'h26C5: d <= 8'hC0; 15'h26C6: d <= 8'hC0; 15'h26C7: d <= 8'hC0;
                15'h26C8: d <= 8'hC0; 15'h26C9: d <= 8'hC0; 15'h26CA: d <= 8'hC0; 15'h26CB: d <= 8'hC0;
                15'h26CC: d <= 8'hC0; 15'h26CD: d <= 8'hC0; 15'h26CE: d <= 8'hC0; 15'h26CF: d <= 8'hC0;
                15'h26D0: d <= 8'hC0; 15'h26D1: d <= 8'hC0; 15'h26D2: d <= 8'hC0; 15'h26D3: d <= 8'hC0;
                15'h26D4: d <= 8'hC0; 15'h26D5: d <= 8'hC0; 15'h26D6: d <= 8'hC0; 15'h26D7: d <= 8'hC0;
                15'h26D8: d <= 8'hC0; 15'h26D9: d <= 8'hC0; 15'h26DA: d <= 8'hC0; 15'h26DB: d <= 8'hC0;
                15'h26DC: d <= 8'hC0; 15'h26DD: d <= 8'hC0; 15'h26DE: d <= 8'hC0; 15'h26DF: d <= 8'hC0;
                15'h26E0: d <= 8'hC0; 15'h26E1: d <= 8'hC0; 15'h26E2: d <= 8'hC0; 15'h26E3: d <= 8'hC0;
                15'h26E4: d <= 8'hC0; 15'h26E5: d <= 8'hC0; 15'h26E6: d <= 8'hC0; 15'h26E7: d <= 8'hC0;
                15'h26E8: d <= 8'hC0; 15'h26E9: d <= 8'hC0; 15'h26EA: d <= 8'hC0; 15'h26EB: d <= 8'hC0;
                15'h26EC: d <= 8'hC0; 15'h26ED: d <= 8'hC0; 15'h26EE: d <= 8'hC0; 15'h26EF: d <= 8'hC0;
                15'h26F0: d <= 8'hC0; 15'h26F1: d <= 8'hC0; 15'h26F2: d <= 8'hC0; 15'h26F3: d <= 8'hC0;
                15'h26F4: d <= 8'hC0; 15'h26F5: d <= 8'hC0; 15'h26F6: d <= 8'hC0; 15'h26F7: d <= 8'hC0;
                15'h26F8: d <= 8'hC0; 15'h26F9: d <= 8'hC0; 15'h26FA: d <= 8'hC0; 15'h26FB: d <= 8'hC0;
                15'h26FC: d <= 8'hC0; 15'h26FD: d <= 8'hC0; 15'h26FE: d <= 8'hC0; 15'h26FF: d <= 8'hC0;
                15'h2700: d <= 8'hC0; 15'h2701: d <= 8'hC0; 15'h2702: d <= 8'hC0; 15'h2703: d <= 8'hC0;
                15'h2704: d <= 8'hC0; 15'h2705: d <= 8'hC0; 15'h2706: d <= 8'hC0; 15'h2707: d <= 8'hC0;
                15'h2708: d <= 8'hC0; 15'h2709: d <= 8'hC0; 15'h270A: d <= 8'hC0; 15'h270B: d <= 8'hC0;
                15'h270C: d <= 8'hC0; 15'h270D: d <= 8'hC0; 15'h270E: d <= 8'hC0; 15'h270F: d <= 8'hC0;
                15'h2710: d <= 8'hC0; 15'h2711: d <= 8'hC0; 15'h2712: d <= 8'hC0; 15'h2713: d <= 8'hC0;
                15'h2714: d <= 8'hC0; 15'h2715: d <= 8'hC0; 15'h2716: d <= 8'hC0; 15'h2717: d <= 8'hC0;
                15'h2718: d <= 8'hC0; 15'h2719: d <= 8'hC0; 15'h271A: d <= 8'hC0; 15'h271B: d <= 8'hC0;
                15'h271C: d <= 8'hC0; 15'h271D: d <= 8'hC0; 15'h271E: d <= 8'hC0; 15'h271F: d <= 8'hC0;
                15'h2720: d <= 8'hC0; 15'h2721: d <= 8'hC0; 15'h2722: d <= 8'hC0; 15'h2723: d <= 8'hC0;
                15'h2724: d <= 8'hC0; 15'h2725: d <= 8'hC0; 15'h2726: d <= 8'hC0; 15'h2727: d <= 8'hC0;
                15'h2728: d <= 8'hC0; 15'h2729: d <= 8'hC0; 15'h272A: d <= 8'hC0; 15'h272B: d <= 8'hC0;
                15'h272C: d <= 8'hC0; 15'h272D: d <= 8'hC0; 15'h272E: d <= 8'hC0; 15'h272F: d <= 8'hC0;
                15'h2730: d <= 8'hC0; 15'h2731: d <= 8'hC0; 15'h2732: d <= 8'hC0; 15'h2733: d <= 8'hC0;
                15'h2734: d <= 8'hC0; 15'h2735: d <= 8'hC0; 15'h2736: d <= 8'hC0; 15'h2737: d <= 8'hC0;
                15'h2738: d <= 8'hC0; 15'h2739: d <= 8'hC0; 15'h273A: d <= 8'hC0; 15'h273B: d <= 8'hC0;
                15'h273C: d <= 8'hC0; 15'h273D: d <= 8'hC0; 15'h273E: d <= 8'hC0; 15'h273F: d <= 8'hC0;
                15'h2740: d <= 8'hC0; 15'h2741: d <= 8'hC0; 15'h2742: d <= 8'hC0; 15'h2743: d <= 8'hC0;
                15'h2744: d <= 8'hC0; 15'h2745: d <= 8'hC0; 15'h2746: d <= 8'hC0; 15'h2747: d <= 8'hC0;
                15'h2748: d <= 8'hC0; 15'h2749: d <= 8'hC0; 15'h274A: d <= 8'hC0; 15'h274B: d <= 8'hC0;
                15'h274C: d <= 8'hC0; 15'h274D: d <= 8'hC0; 15'h274E: d <= 8'hC0; 15'h274F: d <= 8'hC0;
                15'h2750: d <= 8'hC0; 15'h2751: d <= 8'hC0; 15'h2752: d <= 8'hC0; 15'h2753: d <= 8'hC0;
                15'h2754: d <= 8'hC0; 15'h2755: d <= 8'hC0; 15'h2756: d <= 8'hC0; 15'h2757: d <= 8'hC0;
                15'h2758: d <= 8'hC0; 15'h2759: d <= 8'hC0; 15'h275A: d <= 8'hC0; 15'h275B: d <= 8'hC0;
                15'h275C: d <= 8'hC0; 15'h275D: d <= 8'hC0; 15'h275E: d <= 8'hC0; 15'h275F: d <= 8'hC0;
                15'h2760: d <= 8'hC0; 15'h2761: d <= 8'hC0; 15'h2762: d <= 8'hC0; 15'h2763: d <= 8'hC0;
                15'h2764: d <= 8'hC0; 15'h2765: d <= 8'hC0; 15'h2766: d <= 8'hC0; 15'h2767: d <= 8'hC0;
                15'h2768: d <= 8'hC0; 15'h2769: d <= 8'hC0; 15'h276A: d <= 8'hC0; 15'h276B: d <= 8'hC0;
                15'h276C: d <= 8'hC0; 15'h276D: d <= 8'hC0; 15'h276E: d <= 8'hC0; 15'h276F: d <= 8'hC0;
                15'h2770: d <= 8'hC0; 15'h2771: d <= 8'hC0; 15'h2772: d <= 8'hC0; 15'h2773: d <= 8'hC0;
                15'h2774: d <= 8'hC0; 15'h2775: d <= 8'hC0; 15'h2776: d <= 8'hC0; 15'h2777: d <= 8'hC0;
                15'h2778: d <= 8'hC0; 15'h2779: d <= 8'hC0; 15'h277A: d <= 8'hC0; 15'h277B: d <= 8'hC0;
                15'h277C: d <= 8'hC0; 15'h277D: d <= 8'hC0; 15'h277E: d <= 8'hC0; 15'h277F: d <= 8'hC0;
                15'h2780: d <= 8'hC0; 15'h2781: d <= 8'hC0; 15'h2782: d <= 8'hC0; 15'h2783: d <= 8'hC0;
                15'h2784: d <= 8'hC0; 15'h2785: d <= 8'hC0; 15'h2786: d <= 8'hC0; 15'h2787: d <= 8'hC0;
                15'h2788: d <= 8'hC0; 15'h2789: d <= 8'hC0; 15'h278A: d <= 8'hC0; 15'h278B: d <= 8'hC0;
                15'h278C: d <= 8'hC0; 15'h278D: d <= 8'hC0; 15'h278E: d <= 8'hC0; 15'h278F: d <= 8'hC0;
                15'h2790: d <= 8'hC0; 15'h2791: d <= 8'hC0; 15'h2792: d <= 8'hC0; 15'h2793: d <= 8'hC0;
                15'h2794: d <= 8'hC0; 15'h2795: d <= 8'hC0; 15'h2796: d <= 8'hC0; 15'h2797: d <= 8'hC0;
                15'h2798: d <= 8'hC0; 15'h2799: d <= 8'hC0; 15'h279A: d <= 8'hC0; 15'h279B: d <= 8'hC0;
                15'h279C: d <= 8'hC0; 15'h279D: d <= 8'hC0; 15'h279E: d <= 8'hC0; 15'h279F: d <= 8'hC0;
                15'h27A0: d <= 8'hC0; 15'h27A1: d <= 8'hC0; 15'h27A2: d <= 8'hC0; 15'h27A3: d <= 8'hC0;
                15'h27A4: d <= 8'hC0; 15'h27A5: d <= 8'hC0; 15'h27A6: d <= 8'hC0; 15'h27A7: d <= 8'hC0;
                15'h27A8: d <= 8'hC0; 15'h27A9: d <= 8'hC0; 15'h27AA: d <= 8'hC0; 15'h27AB: d <= 8'hC0;
                15'h27AC: d <= 8'hC0; 15'h27AD: d <= 8'hC0; 15'h27AE: d <= 8'hC0; 15'h27AF: d <= 8'hC0;
                15'h27B0: d <= 8'hC0; 15'h27B1: d <= 8'hC0; 15'h27B2: d <= 8'hC0; 15'h27B3: d <= 8'hC0;
                15'h27B4: d <= 8'hC0; 15'h27B5: d <= 8'hC0; 15'h27B6: d <= 8'hC0; 15'h27B7: d <= 8'hC0;
                15'h27B8: d <= 8'hC0; 15'h27B9: d <= 8'hC0; 15'h27BA: d <= 8'hC0; 15'h27BB: d <= 8'hC0;
                15'h27BC: d <= 8'hC0; 15'h27BD: d <= 8'hC0; 15'h27BE: d <= 8'hC0; 15'h27BF: d <= 8'hC0;
                15'h27C0: d <= 8'hC0; 15'h27C1: d <= 8'hC0; 15'h27C2: d <= 8'hC0; 15'h27C3: d <= 8'hC0;
                15'h27C4: d <= 8'hC0; 15'h27C5: d <= 8'hC0; 15'h27C6: d <= 8'hC0; 15'h27C7: d <= 8'hC0;
                15'h27C8: d <= 8'hC0; 15'h27C9: d <= 8'hC0; 15'h27CA: d <= 8'hC0; 15'h27CB: d <= 8'hC0;
                15'h27CC: d <= 8'hC0; 15'h27CD: d <= 8'hC0; 15'h27CE: d <= 8'hC0; 15'h27CF: d <= 8'hC0;
                15'h27D0: d <= 8'hC0; 15'h27D1: d <= 8'hC0; 15'h27D2: d <= 8'hC0; 15'h27D3: d <= 8'hC0;
                15'h27D4: d <= 8'hC0; 15'h27D5: d <= 8'hC0; 15'h27D6: d <= 8'hC0; 15'h27D7: d <= 8'hC0;
                15'h27D8: d <= 8'hC0; 15'h27D9: d <= 8'hC0; 15'h27DA: d <= 8'hC0; 15'h27DB: d <= 8'hC0;
                15'h27DC: d <= 8'hC0; 15'h27DD: d <= 8'hC0; 15'h27DE: d <= 8'hC0; 15'h27DF: d <= 8'hC0;
                15'h27E0: d <= 8'hC0; 15'h27E1: d <= 8'hC0; 15'h27E2: d <= 8'hC0; 15'h27E3: d <= 8'hC0;
                15'h27E4: d <= 8'hC0; 15'h27E5: d <= 8'hC0; 15'h27E6: d <= 8'hC0; 15'h27E7: d <= 8'hC0;
                15'h27E8: d <= 8'hC0; 15'h27E9: d <= 8'hC0; 15'h27EA: d <= 8'hC0; 15'h27EB: d <= 8'hC0;
                15'h27EC: d <= 8'hC0; 15'h27ED: d <= 8'hC0; 15'h27EE: d <= 8'hC0; 15'h27EF: d <= 8'hC0;
                15'h27F0: d <= 8'hC0; 15'h27F1: d <= 8'hC0; 15'h27F2: d <= 8'hC0; 15'h27F3: d <= 8'hC0;
                15'h27F4: d <= 8'hC0; 15'h27F5: d <= 8'hC0; 15'h27F6: d <= 8'hC0; 15'h27F7: d <= 8'hC0;
                15'h27F8: d <= 8'hC0; 15'h27F9: d <= 8'hC0; 15'h27FA: d <= 8'hC0; 15'h27FB: d <= 8'hC0;
                15'h27FC: d <= 8'hC0; 15'h27FD: d <= 8'hC0; 15'h27FE: d <= 8'hC0; 15'h27FF: d <= 8'hC0;
                15'h2800: d <= 8'hC0; 15'h2801: d <= 8'hC0; 15'h2802: d <= 8'hC0; 15'h2803: d <= 8'hC0;
                15'h2804: d <= 8'hC0; 15'h2805: d <= 8'hC0; 15'h2806: d <= 8'hC0; 15'h2807: d <= 8'hC0;
                15'h2808: d <= 8'hC0; 15'h2809: d <= 8'hC0; 15'h280A: d <= 8'hC0; 15'h280B: d <= 8'hC0;
                15'h280C: d <= 8'hC0; 15'h280D: d <= 8'hC0; 15'h280E: d <= 8'hC0; 15'h280F: d <= 8'hC0;
                15'h2810: d <= 8'hC0; 15'h2811: d <= 8'hC0; 15'h2812: d <= 8'hC0; 15'h2813: d <= 8'hC0;
                15'h2814: d <= 8'hC0; 15'h2815: d <= 8'hC0; 15'h2816: d <= 8'hC0; 15'h2817: d <= 8'hC0;
                15'h2818: d <= 8'hC0; 15'h2819: d <= 8'hC0; 15'h281A: d <= 8'hC0; 15'h281B: d <= 8'hC0;
                15'h281C: d <= 8'hC0; 15'h281D: d <= 8'hC0; 15'h281E: d <= 8'hC0; 15'h281F: d <= 8'hC0;
                15'h2820: d <= 8'hC0; 15'h2821: d <= 8'hC0; 15'h2822: d <= 8'hC0; 15'h2823: d <= 8'hC0;
                15'h2824: d <= 8'hC0; 15'h2825: d <= 8'hC0; 15'h2826: d <= 8'hC0; 15'h2827: d <= 8'hC0;
                15'h2828: d <= 8'hC0; 15'h2829: d <= 8'hC0; 15'h282A: d <= 8'hC0; 15'h282B: d <= 8'hC0;
                15'h282C: d <= 8'hC0; 15'h282D: d <= 8'hC0; 15'h282E: d <= 8'hC0; 15'h282F: d <= 8'hC0;
                15'h2830: d <= 8'hC0; 15'h2831: d <= 8'hC0; 15'h2832: d <= 8'hC0; 15'h2833: d <= 8'hC0;
                15'h2834: d <= 8'hC0; 15'h2835: d <= 8'hC0; 15'h2836: d <= 8'hC0; 15'h2837: d <= 8'hC0;
                15'h2838: d <= 8'hC0; 15'h2839: d <= 8'hC0; 15'h283A: d <= 8'hC0; 15'h283B: d <= 8'hC0;
                15'h283C: d <= 8'hC0; 15'h283D: d <= 8'hC0; 15'h283E: d <= 8'hC0; 15'h283F: d <= 8'hC0;
                15'h2840: d <= 8'hC0; 15'h2841: d <= 8'hC0; 15'h2842: d <= 8'hC0; 15'h2843: d <= 8'hC0;
                15'h2844: d <= 8'hC0; 15'h2845: d <= 8'hC0; 15'h2846: d <= 8'hC0; 15'h2847: d <= 8'hC0;
                15'h2848: d <= 8'hC0; 15'h2849: d <= 8'hC0; 15'h284A: d <= 8'hC0; 15'h284B: d <= 8'hC0;
                15'h284C: d <= 8'hC0; 15'h284D: d <= 8'hC0; 15'h284E: d <= 8'hC0; 15'h284F: d <= 8'hC0;
                15'h2850: d <= 8'hC0; 15'h2851: d <= 8'hC0; 15'h2852: d <= 8'hC0; 15'h2853: d <= 8'hC0;
                15'h2854: d <= 8'hC0; 15'h2855: d <= 8'hC0; 15'h2856: d <= 8'hC0; 15'h2857: d <= 8'hC0;
                15'h2858: d <= 8'hC0; 15'h2859: d <= 8'hC0; 15'h285A: d <= 8'hC0; 15'h285B: d <= 8'hC0;
                15'h285C: d <= 8'hC0; 15'h285D: d <= 8'hC0; 15'h285E: d <= 8'hC0; 15'h285F: d <= 8'hC0;
                15'h2860: d <= 8'hC0; 15'h2861: d <= 8'hC0; 15'h2862: d <= 8'hC0; 15'h2863: d <= 8'hC0;
                15'h2864: d <= 8'hC0; 15'h2865: d <= 8'hC0; 15'h2866: d <= 8'hC0; 15'h2867: d <= 8'hC0;
                15'h2868: d <= 8'hC0; 15'h2869: d <= 8'hC0; 15'h286A: d <= 8'hC0; 15'h286B: d <= 8'hC0;
                15'h286C: d <= 8'hC0; 15'h286D: d <= 8'hC0; 15'h286E: d <= 8'hC0; 15'h286F: d <= 8'hC0;
                15'h2870: d <= 8'hC0; 15'h2871: d <= 8'hC0; 15'h2872: d <= 8'hC0; 15'h2873: d <= 8'hC0;
                15'h2874: d <= 8'hC0; 15'h2875: d <= 8'hC0; 15'h2876: d <= 8'hC0; 15'h2877: d <= 8'hC0;
                15'h2878: d <= 8'hC0; 15'h2879: d <= 8'hC0; 15'h287A: d <= 8'hC0; 15'h287B: d <= 8'hC0;
                15'h287C: d <= 8'hC0; 15'h287D: d <= 8'hC0; 15'h287E: d <= 8'hC0; 15'h287F: d <= 8'hC0;
                15'h2880: d <= 8'hC0; 15'h2881: d <= 8'hC0; 15'h2882: d <= 8'hC0; 15'h2883: d <= 8'hC0;
                15'h2884: d <= 8'hC0; 15'h2885: d <= 8'hC0; 15'h2886: d <= 8'hC0; 15'h2887: d <= 8'hC0;
                15'h2888: d <= 8'hC0; 15'h2889: d <= 8'hC0; 15'h288A: d <= 8'hC0; 15'h288B: d <= 8'hC0;
                15'h288C: d <= 8'hC0; 15'h288D: d <= 8'hC0; 15'h288E: d <= 8'hC0; 15'h288F: d <= 8'hC0;
                15'h2890: d <= 8'hC0; 15'h2891: d <= 8'hC0; 15'h2892: d <= 8'hC0; 15'h2893: d <= 8'hC0;
                15'h2894: d <= 8'hC0; 15'h2895: d <= 8'hC0; 15'h2896: d <= 8'hC0; 15'h2897: d <= 8'hC0;
                15'h2898: d <= 8'hC0; 15'h2899: d <= 8'hC0; 15'h289A: d <= 8'hC0; 15'h289B: d <= 8'hC0;
                15'h289C: d <= 8'hC0; 15'h289D: d <= 8'hC0; 15'h289E: d <= 8'hC0; 15'h289F: d <= 8'hC0;
                15'h28A0: d <= 8'hC0; 15'h28A1: d <= 8'hC0; 15'h28A2: d <= 8'hC0; 15'h28A3: d <= 8'hC0;
                15'h28A4: d <= 8'hC0; 15'h28A5: d <= 8'hC0; 15'h28A6: d <= 8'hC0; 15'h28A7: d <= 8'hC0;
                15'h28A8: d <= 8'hC0; 15'h28A9: d <= 8'hC0; 15'h28AA: d <= 8'hC0; 15'h28AB: d <= 8'hC0;
                15'h28AC: d <= 8'hC0; 15'h28AD: d <= 8'hC0; 15'h28AE: d <= 8'hC0; 15'h28AF: d <= 8'hC0;
                15'h28B0: d <= 8'hC0; 15'h28B1: d <= 8'hC0; 15'h28B2: d <= 8'hC0; 15'h28B3: d <= 8'hC0;
                15'h28B4: d <= 8'hC0; 15'h28B5: d <= 8'hC0; 15'h28B6: d <= 8'hC0; 15'h28B7: d <= 8'hC0;
                15'h28B8: d <= 8'hC0; 15'h28B9: d <= 8'hC0; 15'h28BA: d <= 8'hC0; 15'h28BB: d <= 8'hC0;
                15'h28BC: d <= 8'hC0; 15'h28BD: d <= 8'hC0; 15'h28BE: d <= 8'hC0; 15'h28BF: d <= 8'hC0;
                15'h28C0: d <= 8'hC0; 15'h28C1: d <= 8'hC0; 15'h28C2: d <= 8'hC0; 15'h28C3: d <= 8'hC0;
                15'h28C4: d <= 8'hC0; 15'h28C5: d <= 8'hC0; 15'h28C6: d <= 8'hC0; 15'h28C7: d <= 8'hC0;
                15'h28C8: d <= 8'hC0; 15'h28C9: d <= 8'hC0; 15'h28CA: d <= 8'hC0; 15'h28CB: d <= 8'hC0;
                15'h28CC: d <= 8'hC0; 15'h28CD: d <= 8'hC0; 15'h28CE: d <= 8'hC0; 15'h28CF: d <= 8'hC0;
                15'h28D0: d <= 8'hC0; 15'h28D1: d <= 8'hC0; 15'h28D2: d <= 8'hC0; 15'h28D3: d <= 8'hC0;
                15'h28D4: d <= 8'hC0; 15'h28D5: d <= 8'hC0; 15'h28D6: d <= 8'hC0; 15'h28D7: d <= 8'hC0;
                15'h28D8: d <= 8'hC0; 15'h28D9: d <= 8'hC0; 15'h28DA: d <= 8'hC0; 15'h28DB: d <= 8'hC0;
                15'h28DC: d <= 8'hC0; 15'h28DD: d <= 8'hC0; 15'h28DE: d <= 8'hC0; 15'h28DF: d <= 8'hC0;
                15'h28E0: d <= 8'hC0; 15'h28E1: d <= 8'hC0; 15'h28E2: d <= 8'hC0; 15'h28E3: d <= 8'hC0;
                15'h28E4: d <= 8'hC0; 15'h28E5: d <= 8'hC0; 15'h28E6: d <= 8'hC0; 15'h28E7: d <= 8'hC0;
                15'h28E8: d <= 8'hC0; 15'h28E9: d <= 8'hC0; 15'h28EA: d <= 8'hC0; 15'h28EB: d <= 8'hC0;
                15'h28EC: d <= 8'hC0; 15'h28ED: d <= 8'hC0; 15'h28EE: d <= 8'hC0; 15'h28EF: d <= 8'hC0;
                15'h28F0: d <= 8'hC0; 15'h28F1: d <= 8'hC0; 15'h28F2: d <= 8'hC0; 15'h28F3: d <= 8'hC0;
                15'h28F4: d <= 8'hC0; 15'h28F5: d <= 8'hC0; 15'h28F6: d <= 8'hC0; 15'h28F7: d <= 8'hC0;
                15'h28F8: d <= 8'hC0; 15'h28F9: d <= 8'hC0; 15'h28FA: d <= 8'hC0; 15'h28FB: d <= 8'hC0;
                15'h28FC: d <= 8'hC0; 15'h28FD: d <= 8'hC0; 15'h28FE: d <= 8'hC0; 15'h28FF: d <= 8'hC0;
                15'h2900: d <= 8'hC0; 15'h2901: d <= 8'hC0; 15'h2902: d <= 8'hC0; 15'h2903: d <= 8'hC0;
                15'h2904: d <= 8'hC0; 15'h2905: d <= 8'hC0; 15'h2906: d <= 8'hC0; 15'h2907: d <= 8'hC0;
                15'h2908: d <= 8'hC0; 15'h2909: d <= 8'hC0; 15'h290A: d <= 8'hC0; 15'h290B: d <= 8'hC0;
                15'h290C: d <= 8'hC0; 15'h290D: d <= 8'hC0; 15'h290E: d <= 8'hC0; 15'h290F: d <= 8'hC0;
                15'h2910: d <= 8'hC0; 15'h2911: d <= 8'hC0; 15'h2912: d <= 8'hC0; 15'h2913: d <= 8'hC0;
                15'h2914: d <= 8'hC0; 15'h2915: d <= 8'hC0; 15'h2916: d <= 8'hC0; 15'h2917: d <= 8'hC0;
                15'h2918: d <= 8'hC0; 15'h2919: d <= 8'hC0; 15'h291A: d <= 8'hC0; 15'h291B: d <= 8'hC0;
                15'h291C: d <= 8'hC0; 15'h291D: d <= 8'hC0; 15'h291E: d <= 8'hC0; 15'h291F: d <= 8'hC0;
                15'h2920: d <= 8'hC0; 15'h2921: d <= 8'hC0; 15'h2922: d <= 8'hC0; 15'h2923: d <= 8'hC0;
                15'h2924: d <= 8'hC0; 15'h2925: d <= 8'hC0; 15'h2926: d <= 8'hC0; 15'h2927: d <= 8'hC0;
                15'h2928: d <= 8'hC0; 15'h2929: d <= 8'hC0; 15'h292A: d <= 8'hC0; 15'h292B: d <= 8'hC0;
                15'h292C: d <= 8'hC0; 15'h292D: d <= 8'hC0; 15'h292E: d <= 8'hC0; 15'h292F: d <= 8'hC0;
                15'h2930: d <= 8'hC0; 15'h2931: d <= 8'hC0; 15'h2932: d <= 8'hC0; 15'h2933: d <= 8'hC0;
                15'h2934: d <= 8'hC0; 15'h2935: d <= 8'hC0; 15'h2936: d <= 8'hC0; 15'h2937: d <= 8'hC0;
                15'h2938: d <= 8'hC0; 15'h2939: d <= 8'hC0; 15'h293A: d <= 8'hC0; 15'h293B: d <= 8'hC0;
                15'h293C: d <= 8'hC0; 15'h293D: d <= 8'hC0; 15'h293E: d <= 8'hC0; 15'h293F: d <= 8'hC0;
                15'h2940: d <= 8'hC0; 15'h2941: d <= 8'hC0; 15'h2942: d <= 8'hC0; 15'h2943: d <= 8'hC0;
                15'h2944: d <= 8'hC0; 15'h2945: d <= 8'hC0; 15'h2946: d <= 8'hC0; 15'h2947: d <= 8'hC0;
                15'h2948: d <= 8'hC0; 15'h2949: d <= 8'hC0; 15'h294A: d <= 8'hC0; 15'h294B: d <= 8'hC0;
                15'h294C: d <= 8'hC0; 15'h294D: d <= 8'hC0; 15'h294E: d <= 8'hC0; 15'h294F: d <= 8'hC0;
                15'h2950: d <= 8'hC0; 15'h2951: d <= 8'hC0; 15'h2952: d <= 8'hC0; 15'h2953: d <= 8'hC0;
                15'h2954: d <= 8'hC0; 15'h2955: d <= 8'hC0; 15'h2956: d <= 8'hC0; 15'h2957: d <= 8'hC0;
                15'h2958: d <= 8'hC0; 15'h2959: d <= 8'hC0; 15'h295A: d <= 8'hC0; 15'h295B: d <= 8'hC0;
                15'h295C: d <= 8'hC0; 15'h295D: d <= 8'hC0; 15'h295E: d <= 8'hC0; 15'h295F: d <= 8'hC0;
                15'h2960: d <= 8'hC0; 15'h2961: d <= 8'hC0; 15'h2962: d <= 8'hC0; 15'h2963: d <= 8'hC0;
                15'h2964: d <= 8'hC0; 15'h2965: d <= 8'hC0; 15'h2966: d <= 8'hC0; 15'h2967: d <= 8'hC0;
                15'h2968: d <= 8'hC0; 15'h2969: d <= 8'hC0; 15'h296A: d <= 8'hC0; 15'h296B: d <= 8'hC0;
                15'h296C: d <= 8'hC0; 15'h296D: d <= 8'hC0; 15'h296E: d <= 8'hC0; 15'h296F: d <= 8'hC0;
                15'h2970: d <= 8'hC0; 15'h2971: d <= 8'hC0; 15'h2972: d <= 8'hC0; 15'h2973: d <= 8'hC0;
                15'h2974: d <= 8'hC0; 15'h2975: d <= 8'hC0; 15'h2976: d <= 8'hC0; 15'h2977: d <= 8'hC0;
                15'h2978: d <= 8'hC0; 15'h2979: d <= 8'hC0; 15'h297A: d <= 8'hC0; 15'h297B: d <= 8'hC0;
                15'h297C: d <= 8'hC0; 15'h297D: d <= 8'hC0; 15'h297E: d <= 8'hC0; 15'h297F: d <= 8'hC0;
                15'h2980: d <= 8'hC0; 15'h2981: d <= 8'hC0; 15'h2982: d <= 8'hC0; 15'h2983: d <= 8'hC0;
                15'h2984: d <= 8'hC0; 15'h2985: d <= 8'hC0; 15'h2986: d <= 8'hC0; 15'h2987: d <= 8'hC0;
                15'h2988: d <= 8'hC0; 15'h2989: d <= 8'hC0; 15'h298A: d <= 8'hC0; 15'h298B: d <= 8'hC0;
                15'h298C: d <= 8'hC0; 15'h298D: d <= 8'hC0; 15'h298E: d <= 8'hC0; 15'h298F: d <= 8'hC0;
                15'h2990: d <= 8'hC0; 15'h2991: d <= 8'hC0; 15'h2992: d <= 8'hC0; 15'h2993: d <= 8'hC0;
                15'h2994: d <= 8'hC0; 15'h2995: d <= 8'hC0; 15'h2996: d <= 8'hC0; 15'h2997: d <= 8'hC0;
                15'h2998: d <= 8'hC0; 15'h2999: d <= 8'hC0; 15'h299A: d <= 8'hC0; 15'h299B: d <= 8'hC0;
                15'h299C: d <= 8'hC0; 15'h299D: d <= 8'hC0; 15'h299E: d <= 8'hC0; 15'h299F: d <= 8'hC0;
                15'h29A0: d <= 8'hC0; 15'h29A1: d <= 8'hC0; 15'h29A2: d <= 8'hC0; 15'h29A3: d <= 8'hC0;
                15'h29A4: d <= 8'hC0; 15'h29A5: d <= 8'hC0; 15'h29A6: d <= 8'hC0; 15'h29A7: d <= 8'hC0;
                15'h29A8: d <= 8'hC0; 15'h29A9: d <= 8'hC0; 15'h29AA: d <= 8'hC0; 15'h29AB: d <= 8'hC0;
                15'h29AC: d <= 8'hC0; 15'h29AD: d <= 8'hC0; 15'h29AE: d <= 8'hC0; 15'h29AF: d <= 8'hC0;
                15'h29B0: d <= 8'hC0; 15'h29B1: d <= 8'hC0; 15'h29B2: d <= 8'hC0; 15'h29B3: d <= 8'hC0;
                15'h29B4: d <= 8'hC0; 15'h29B5: d <= 8'hC0; 15'h29B6: d <= 8'hC0; 15'h29B7: d <= 8'hC0;
                15'h29B8: d <= 8'hC0; 15'h29B9: d <= 8'hC0; 15'h29BA: d <= 8'hC0; 15'h29BB: d <= 8'hC0;
                15'h29BC: d <= 8'hC0; 15'h29BD: d <= 8'hC0; 15'h29BE: d <= 8'hC0; 15'h29BF: d <= 8'hC0;
                15'h29C0: d <= 8'hC0; 15'h29C1: d <= 8'hC0; 15'h29C2: d <= 8'hC0; 15'h29C3: d <= 8'hC0;
                15'h29C4: d <= 8'hC0; 15'h29C5: d <= 8'hC0; 15'h29C6: d <= 8'hC0; 15'h29C7: d <= 8'hC0;
                15'h29C8: d <= 8'hC0; 15'h29C9: d <= 8'hC0; 15'h29CA: d <= 8'hC0; 15'h29CB: d <= 8'hC0;
                15'h29CC: d <= 8'hC0; 15'h29CD: d <= 8'hC0; 15'h29CE: d <= 8'hC0; 15'h29CF: d <= 8'hC0;
                15'h29D0: d <= 8'hC0; 15'h29D1: d <= 8'hC0; 15'h29D2: d <= 8'hC0; 15'h29D3: d <= 8'hC0;
                15'h29D4: d <= 8'hC0; 15'h29D5: d <= 8'hC0; 15'h29D6: d <= 8'hC0; 15'h29D7: d <= 8'hC0;
                15'h29D8: d <= 8'hC0; 15'h29D9: d <= 8'hC0; 15'h29DA: d <= 8'hC0; 15'h29DB: d <= 8'hC0;
                15'h29DC: d <= 8'hC0; 15'h29DD: d <= 8'hC0; 15'h29DE: d <= 8'hC0; 15'h29DF: d <= 8'hC0;
                15'h29E0: d <= 8'hC0; 15'h29E1: d <= 8'hC0; 15'h29E2: d <= 8'hC0; 15'h29E3: d <= 8'hC0;
                15'h29E4: d <= 8'hC0; 15'h29E5: d <= 8'hC0; 15'h29E6: d <= 8'hC0; 15'h29E7: d <= 8'hC0;
                15'h29E8: d <= 8'hC0; 15'h29E9: d <= 8'hC0; 15'h29EA: d <= 8'hC0; 15'h29EB: d <= 8'hC0;
                15'h29EC: d <= 8'hC0; 15'h29ED: d <= 8'hC0; 15'h29EE: d <= 8'hC0; 15'h29EF: d <= 8'hC0;
                15'h29F0: d <= 8'hC0; 15'h29F1: d <= 8'hC0; 15'h29F2: d <= 8'hC0; 15'h29F3: d <= 8'hC0;
                15'h29F4: d <= 8'hC0; 15'h29F5: d <= 8'hC0; 15'h29F6: d <= 8'hC0; 15'h29F7: d <= 8'hC0;
                15'h29F8: d <= 8'hC0; 15'h29F9: d <= 8'hC0; 15'h29FA: d <= 8'hC0; 15'h29FB: d <= 8'hC0;
                15'h29FC: d <= 8'hC0; 15'h29FD: d <= 8'hC0; 15'h29FE: d <= 8'hC0; 15'h29FF: d <= 8'hC0;
                15'h2A00: d <= 8'hC0; 15'h2A01: d <= 8'hC0; 15'h2A02: d <= 8'hC0; 15'h2A03: d <= 8'hC0;
                15'h2A04: d <= 8'hC0; 15'h2A05: d <= 8'hC0; 15'h2A06: d <= 8'hC0; 15'h2A07: d <= 8'hC0;
                15'h2A08: d <= 8'hC0; 15'h2A09: d <= 8'hC0; 15'h2A0A: d <= 8'hC0; 15'h2A0B: d <= 8'hC0;
                15'h2A0C: d <= 8'hC0; 15'h2A0D: d <= 8'hC0; 15'h2A0E: d <= 8'hC0; 15'h2A0F: d <= 8'hC0;
                15'h2A10: d <= 8'hC0; 15'h2A11: d <= 8'hC0; 15'h2A12: d <= 8'hC0; 15'h2A13: d <= 8'hC0;
                15'h2A14: d <= 8'hC0; 15'h2A15: d <= 8'hC0; 15'h2A16: d <= 8'hC0; 15'h2A17: d <= 8'hC0;
                15'h2A18: d <= 8'hC0; 15'h2A19: d <= 8'hC0; 15'h2A1A: d <= 8'hC0; 15'h2A1B: d <= 8'hC0;
                15'h2A1C: d <= 8'hC0; 15'h2A1D: d <= 8'hC0; 15'h2A1E: d <= 8'hC0; 15'h2A1F: d <= 8'hC0;
                15'h2A20: d <= 8'hC0; 15'h2A21: d <= 8'hC0; 15'h2A22: d <= 8'hC0; 15'h2A23: d <= 8'hC0;
                15'h2A24: d <= 8'hC0; 15'h2A25: d <= 8'hC0; 15'h2A26: d <= 8'hC0; 15'h2A27: d <= 8'hC0;
                15'h2A28: d <= 8'hC0; 15'h2A29: d <= 8'hC0; 15'h2A2A: d <= 8'hC0; 15'h2A2B: d <= 8'hC0;
                15'h2A2C: d <= 8'hC0; 15'h2A2D: d <= 8'hC0; 15'h2A2E: d <= 8'hC0; 15'h2A2F: d <= 8'hC0;
                15'h2A30: d <= 8'hC0; 15'h2A31: d <= 8'hC0; 15'h2A32: d <= 8'hC0; 15'h2A33: d <= 8'hC0;
                15'h2A34: d <= 8'hC0; 15'h2A35: d <= 8'hC0; 15'h2A36: d <= 8'hC0; 15'h2A37: d <= 8'hC0;
                15'h2A38: d <= 8'hC0; 15'h2A39: d <= 8'hC0; 15'h2A3A: d <= 8'hC0; 15'h2A3B: d <= 8'hC0;
                15'h2A3C: d <= 8'hC0; 15'h2A3D: d <= 8'hC0; 15'h2A3E: d <= 8'hC0; 15'h2A3F: d <= 8'hC0;
                15'h2A40: d <= 8'hC0; 15'h2A41: d <= 8'hC0; 15'h2A42: d <= 8'hC0; 15'h2A43: d <= 8'hC0;
                15'h2A44: d <= 8'hC0; 15'h2A45: d <= 8'hC0; 15'h2A46: d <= 8'hC0; 15'h2A47: d <= 8'hC0;
                15'h2A48: d <= 8'hC0; 15'h2A49: d <= 8'hC0; 15'h2A4A: d <= 8'hC0; 15'h2A4B: d <= 8'hC0;
                15'h2A4C: d <= 8'hC0; 15'h2A4D: d <= 8'hC0; 15'h2A4E: d <= 8'hC0; 15'h2A4F: d <= 8'hC0;
                15'h2A50: d <= 8'hC0; 15'h2A51: d <= 8'hC0; 15'h2A52: d <= 8'hC0; 15'h2A53: d <= 8'hC0;
                15'h2A54: d <= 8'hC0; 15'h2A55: d <= 8'hC0; 15'h2A56: d <= 8'hC0; 15'h2A57: d <= 8'hC0;
                15'h2A58: d <= 8'hC0; 15'h2A59: d <= 8'hC0; 15'h2A5A: d <= 8'hC0; 15'h2A5B: d <= 8'hC0;
                15'h2A5C: d <= 8'hC0; 15'h2A5D: d <= 8'hC0; 15'h2A5E: d <= 8'hC0; 15'h2A5F: d <= 8'hC0;
                15'h2A60: d <= 8'hC0; 15'h2A61: d <= 8'hC0; 15'h2A62: d <= 8'hC0; 15'h2A63: d <= 8'hC0;
                15'h2A64: d <= 8'hC0; 15'h2A65: d <= 8'hC0; 15'h2A66: d <= 8'hC0; 15'h2A67: d <= 8'hC0;
                15'h2A68: d <= 8'hC0; 15'h2A69: d <= 8'hC0; 15'h2A6A: d <= 8'hC0; 15'h2A6B: d <= 8'hC0;
                15'h2A6C: d <= 8'hC0; 15'h2A6D: d <= 8'hC0; 15'h2A6E: d <= 8'hC0; 15'h2A6F: d <= 8'hC0;
                15'h2A70: d <= 8'hC0; 15'h2A71: d <= 8'hC0; 15'h2A72: d <= 8'hC0; 15'h2A73: d <= 8'hC0;
                15'h2A74: d <= 8'hC0; 15'h2A75: d <= 8'hC0; 15'h2A76: d <= 8'hC0; 15'h2A77: d <= 8'hC0;
                15'h2A78: d <= 8'hC0; 15'h2A79: d <= 8'hC0; 15'h2A7A: d <= 8'hC0; 15'h2A7B: d <= 8'hC0;
                15'h2A7C: d <= 8'hC0; 15'h2A7D: d <= 8'hC0; 15'h2A7E: d <= 8'hC0; 15'h2A7F: d <= 8'hC0;
                15'h2A80: d <= 8'hC0; 15'h2A81: d <= 8'hC0; 15'h2A82: d <= 8'hC0; 15'h2A83: d <= 8'hC0;
                15'h2A84: d <= 8'hC0; 15'h2A85: d <= 8'hC0; 15'h2A86: d <= 8'hC0; 15'h2A87: d <= 8'hC0;
                15'h2A88: d <= 8'hC0; 15'h2A89: d <= 8'hC0; 15'h2A8A: d <= 8'hC0; 15'h2A8B: d <= 8'hC0;
                15'h2A8C: d <= 8'hC0; 15'h2A8D: d <= 8'hC0; 15'h2A8E: d <= 8'hC0; 15'h2A8F: d <= 8'hC0;
                15'h2A90: d <= 8'hC0; 15'h2A91: d <= 8'hC0; 15'h2A92: d <= 8'hC0; 15'h2A93: d <= 8'hC0;
                15'h2A94: d <= 8'hC0; 15'h2A95: d <= 8'hC0; 15'h2A96: d <= 8'hC0; 15'h2A97: d <= 8'hC0;
                15'h2A98: d <= 8'hC0; 15'h2A99: d <= 8'hC0; 15'h2A9A: d <= 8'hC0; 15'h2A9B: d <= 8'hC0;
                15'h2A9C: d <= 8'hC0; 15'h2A9D: d <= 8'hC0; 15'h2A9E: d <= 8'hC0; 15'h2A9F: d <= 8'hC0;
                15'h2AA0: d <= 8'hC0; 15'h2AA1: d <= 8'hC0; 15'h2AA2: d <= 8'hC0; 15'h2AA3: d <= 8'hC0;
                15'h2AA4: d <= 8'hC0; 15'h2AA5: d <= 8'hC0; 15'h2AA6: d <= 8'hC0; 15'h2AA7: d <= 8'hC0;
                15'h2AA8: d <= 8'hC0; 15'h2AA9: d <= 8'hC0; 15'h2AAA: d <= 8'hC0; 15'h2AAB: d <= 8'hC0;
                15'h2AAC: d <= 8'hC0; 15'h2AAD: d <= 8'hC0; 15'h2AAE: d <= 8'hC0; 15'h2AAF: d <= 8'hC0;
                15'h2AB0: d <= 8'hC0; 15'h2AB1: d <= 8'hC0; 15'h2AB2: d <= 8'hC0; 15'h2AB3: d <= 8'hC0;
                15'h2AB4: d <= 8'hC0; 15'h2AB5: d <= 8'hC0; 15'h2AB6: d <= 8'hC0; 15'h2AB7: d <= 8'hC0;
                15'h2AB8: d <= 8'hC0; 15'h2AB9: d <= 8'hC0; 15'h2ABA: d <= 8'hC0; 15'h2ABB: d <= 8'hC0;
                15'h2ABC: d <= 8'hC0; 15'h2ABD: d <= 8'hC0; 15'h2ABE: d <= 8'hC0; 15'h2ABF: d <= 8'hC0;
                15'h2AC0: d <= 8'hC0; 15'h2AC1: d <= 8'hC0; 15'h2AC2: d <= 8'hC0; 15'h2AC3: d <= 8'hC0;
                15'h2AC4: d <= 8'hC0; 15'h2AC5: d <= 8'hC0; 15'h2AC6: d <= 8'hC0; 15'h2AC7: d <= 8'hC0;
                15'h2AC8: d <= 8'hC0; 15'h2AC9: d <= 8'hC0; 15'h2ACA: d <= 8'hC0; 15'h2ACB: d <= 8'hC0;
                15'h2ACC: d <= 8'hC0; 15'h2ACD: d <= 8'hC0; 15'h2ACE: d <= 8'hC0; 15'h2ACF: d <= 8'hC0;
                15'h2AD0: d <= 8'hC0; 15'h2AD1: d <= 8'hC0; 15'h2AD2: d <= 8'hC0; 15'h2AD3: d <= 8'hC0;
                15'h2AD4: d <= 8'hC0; 15'h2AD5: d <= 8'hC0; 15'h2AD6: d <= 8'hC0; 15'h2AD7: d <= 8'hC0;
                15'h2AD8: d <= 8'hC0; 15'h2AD9: d <= 8'hC0; 15'h2ADA: d <= 8'hC0; 15'h2ADB: d <= 8'hC0;
                15'h2ADC: d <= 8'hC0; 15'h2ADD: d <= 8'hC0; 15'h2ADE: d <= 8'hC0; 15'h2ADF: d <= 8'hC0;
                15'h2AE0: d <= 8'hC0; 15'h2AE1: d <= 8'hC0; 15'h2AE2: d <= 8'hC0; 15'h2AE3: d <= 8'hC0;
                15'h2AE4: d <= 8'hC0; 15'h2AE5: d <= 8'hC0; 15'h2AE6: d <= 8'hC0; 15'h2AE7: d <= 8'hC0;
                15'h2AE8: d <= 8'hC0; 15'h2AE9: d <= 8'hC0; 15'h2AEA: d <= 8'hC0; 15'h2AEB: d <= 8'hC0;
                15'h2AEC: d <= 8'hC0; 15'h2AED: d <= 8'hC0; 15'h2AEE: d <= 8'hC0; 15'h2AEF: d <= 8'hC0;
                15'h2AF0: d <= 8'hC0; 15'h2AF1: d <= 8'hC0; 15'h2AF2: d <= 8'hC0; 15'h2AF3: d <= 8'hC0;
                15'h2AF4: d <= 8'hC0; 15'h2AF5: d <= 8'hC0; 15'h2AF6: d <= 8'hC0; 15'h2AF7: d <= 8'hC0;
                15'h2AF8: d <= 8'hC0; 15'h2AF9: d <= 8'hC0; 15'h2AFA: d <= 8'hC0; 15'h2AFB: d <= 8'hC0;
                15'h2AFC: d <= 8'hC0; 15'h2AFD: d <= 8'hC0; 15'h2AFE: d <= 8'hC0; 15'h2AFF: d <= 8'hC0;
                15'h2B00: d <= 8'hC0; 15'h2B01: d <= 8'hC0; 15'h2B02: d <= 8'hC0; 15'h2B03: d <= 8'hC0;
                15'h2B04: d <= 8'hC0; 15'h2B05: d <= 8'hC0; 15'h2B06: d <= 8'hC0; 15'h2B07: d <= 8'hC0;
                15'h2B08: d <= 8'hC0; 15'h2B09: d <= 8'hC0; 15'h2B0A: d <= 8'hC0; 15'h2B0B: d <= 8'hC0;
                15'h2B0C: d <= 8'hC0; 15'h2B0D: d <= 8'hC0; 15'h2B0E: d <= 8'hC0; 15'h2B0F: d <= 8'hC0;
                15'h2B10: d <= 8'hC0; 15'h2B11: d <= 8'hC0; 15'h2B12: d <= 8'hC0; 15'h2B13: d <= 8'hC0;
                15'h2B14: d <= 8'hC0; 15'h2B15: d <= 8'hC0; 15'h2B16: d <= 8'hC0; 15'h2B17: d <= 8'hC0;
                15'h2B18: d <= 8'hC0; 15'h2B19: d <= 8'hC0; 15'h2B1A: d <= 8'hC0; 15'h2B1B: d <= 8'hC0;
                15'h2B1C: d <= 8'hC0; 15'h2B1D: d <= 8'hC0; 15'h2B1E: d <= 8'hC0; 15'h2B1F: d <= 8'hC0;
                15'h2B20: d <= 8'hC0; 15'h2B21: d <= 8'hC0; 15'h2B22: d <= 8'hC0; 15'h2B23: d <= 8'hC0;
                15'h2B24: d <= 8'hC0; 15'h2B25: d <= 8'hC0; 15'h2B26: d <= 8'hC0; 15'h2B27: d <= 8'hC0;
                15'h2B28: d <= 8'hC0; 15'h2B29: d <= 8'hC0; 15'h2B2A: d <= 8'hC0; 15'h2B2B: d <= 8'hC0;
                15'h2B2C: d <= 8'hC0; 15'h2B2D: d <= 8'hC0; 15'h2B2E: d <= 8'hC0; 15'h2B2F: d <= 8'hC0;
                15'h2B30: d <= 8'hC0; 15'h2B31: d <= 8'hC0; 15'h2B32: d <= 8'hC0; 15'h2B33: d <= 8'hC0;
                15'h2B34: d <= 8'hC0; 15'h2B35: d <= 8'hC0; 15'h2B36: d <= 8'hC0; 15'h2B37: d <= 8'hC0;
                15'h2B38: d <= 8'hC0; 15'h2B39: d <= 8'hC0; 15'h2B3A: d <= 8'hC0; 15'h2B3B: d <= 8'hC0;
                15'h2B3C: d <= 8'hC0; 15'h2B3D: d <= 8'hC0; 15'h2B3E: d <= 8'hC0; 15'h2B3F: d <= 8'hC0;
                15'h2B40: d <= 8'hC0; 15'h2B41: d <= 8'hC0; 15'h2B42: d <= 8'hC0; 15'h2B43: d <= 8'hC0;
                15'h2B44: d <= 8'hC0; 15'h2B45: d <= 8'hC0; 15'h2B46: d <= 8'hC0; 15'h2B47: d <= 8'hC0;
                15'h2B48: d <= 8'hC0; 15'h2B49: d <= 8'hC0; 15'h2B4A: d <= 8'hC0; 15'h2B4B: d <= 8'hC0;
                15'h2B4C: d <= 8'hC0; 15'h2B4D: d <= 8'hC0; 15'h2B4E: d <= 8'hC0; 15'h2B4F: d <= 8'hC0;
                15'h2B50: d <= 8'hC0; 15'h2B51: d <= 8'hC0; 15'h2B52: d <= 8'hC0; 15'h2B53: d <= 8'hC0;
                15'h2B54: d <= 8'hC0; 15'h2B55: d <= 8'hC0; 15'h2B56: d <= 8'hC0; 15'h2B57: d <= 8'hC0;
                15'h2B58: d <= 8'hC0; 15'h2B59: d <= 8'hC0; 15'h2B5A: d <= 8'hC0; 15'h2B5B: d <= 8'hC0;
                15'h2B5C: d <= 8'hC0; 15'h2B5D: d <= 8'hC0; 15'h2B5E: d <= 8'hC0; 15'h2B5F: d <= 8'hC0;
                15'h2B60: d <= 8'hC0; 15'h2B61: d <= 8'hC0; 15'h2B62: d <= 8'hC0; 15'h2B63: d <= 8'hC0;
                15'h2B64: d <= 8'hC0; 15'h2B65: d <= 8'hC0; 15'h2B66: d <= 8'hC0; 15'h2B67: d <= 8'hC0;
                15'h2B68: d <= 8'hC0; 15'h2B69: d <= 8'hC0; 15'h2B6A: d <= 8'hC0; 15'h2B6B: d <= 8'hC0;
                15'h2B6C: d <= 8'hC0; 15'h2B6D: d <= 8'hC0; 15'h2B6E: d <= 8'hC0; 15'h2B6F: d <= 8'hC0;
                15'h2B70: d <= 8'hC0; 15'h2B71: d <= 8'hC0; 15'h2B72: d <= 8'hC0; 15'h2B73: d <= 8'hC0;
                15'h2B74: d <= 8'hC0; 15'h2B75: d <= 8'hC0; 15'h2B76: d <= 8'hC0; 15'h2B77: d <= 8'hC0;
                15'h2B78: d <= 8'hC0; 15'h2B79: d <= 8'hC0; 15'h2B7A: d <= 8'hC0; 15'h2B7B: d <= 8'hC0;
                15'h2B7C: d <= 8'hC0; 15'h2B7D: d <= 8'hC0; 15'h2B7E: d <= 8'hC0; 15'h2B7F: d <= 8'hC0;
                15'h2B80: d <= 8'hC0; 15'h2B81: d <= 8'hC0; 15'h2B82: d <= 8'hC0; 15'h2B83: d <= 8'hC0;
                15'h2B84: d <= 8'hC0; 15'h2B85: d <= 8'hC0; 15'h2B86: d <= 8'hC0; 15'h2B87: d <= 8'hC0;
                15'h2B88: d <= 8'hC0; 15'h2B89: d <= 8'hC0; 15'h2B8A: d <= 8'hC0; 15'h2B8B: d <= 8'hC0;
                15'h2B8C: d <= 8'hC0; 15'h2B8D: d <= 8'hC0; 15'h2B8E: d <= 8'hC0; 15'h2B8F: d <= 8'hC0;
                15'h2B90: d <= 8'hC0; 15'h2B91: d <= 8'hC0; 15'h2B92: d <= 8'hC0; 15'h2B93: d <= 8'hC0;
                15'h2B94: d <= 8'hC0; 15'h2B95: d <= 8'hC0; 15'h2B96: d <= 8'hC0; 15'h2B97: d <= 8'hC0;
                15'h2B98: d <= 8'hC0; 15'h2B99: d <= 8'hC0; 15'h2B9A: d <= 8'hC0; 15'h2B9B: d <= 8'hC0;
                15'h2B9C: d <= 8'hC0; 15'h2B9D: d <= 8'hC0; 15'h2B9E: d <= 8'hC0; 15'h2B9F: d <= 8'hC0;
                15'h2BA0: d <= 8'hC0; 15'h2BA1: d <= 8'hC0; 15'h2BA2: d <= 8'hC0; 15'h2BA3: d <= 8'hC0;
                15'h2BA4: d <= 8'hC0; 15'h2BA5: d <= 8'hC0; 15'h2BA6: d <= 8'hC0; 15'h2BA7: d <= 8'hC0;
                15'h2BA8: d <= 8'hC0; 15'h2BA9: d <= 8'hC0; 15'h2BAA: d <= 8'hC0; 15'h2BAB: d <= 8'hC0;
                15'h2BAC: d <= 8'hC0; 15'h2BAD: d <= 8'hC0; 15'h2BAE: d <= 8'hC0; 15'h2BAF: d <= 8'hC0;
                15'h2BB0: d <= 8'hC0; 15'h2BB1: d <= 8'hC0; 15'h2BB2: d <= 8'hC0; 15'h2BB3: d <= 8'hC0;
                15'h2BB4: d <= 8'hC0; 15'h2BB5: d <= 8'hC0; 15'h2BB6: d <= 8'hC0; 15'h2BB7: d <= 8'hC0;
                15'h2BB8: d <= 8'hC0; 15'h2BB9: d <= 8'hC0; 15'h2BBA: d <= 8'hC0; 15'h2BBB: d <= 8'hC0;
                15'h2BBC: d <= 8'hC0; 15'h2BBD: d <= 8'hC0; 15'h2BBE: d <= 8'hC0; 15'h2BBF: d <= 8'hC0;
                15'h2BC0: d <= 8'hC0; 15'h2BC1: d <= 8'hC0; 15'h2BC2: d <= 8'hC0; 15'h2BC3: d <= 8'hC0;
                15'h2BC4: d <= 8'hC0; 15'h2BC5: d <= 8'hC0; 15'h2BC6: d <= 8'hC0; 15'h2BC7: d <= 8'hC0;
                15'h2BC8: d <= 8'hC0; 15'h2BC9: d <= 8'hC0; 15'h2BCA: d <= 8'hC0; 15'h2BCB: d <= 8'hC0;
                15'h2BCC: d <= 8'hC0; 15'h2BCD: d <= 8'hC0; 15'h2BCE: d <= 8'hC0; 15'h2BCF: d <= 8'hC0;
                15'h2BD0: d <= 8'hC0; 15'h2BD1: d <= 8'hC0; 15'h2BD2: d <= 8'hC0; 15'h2BD3: d <= 8'hC0;
                15'h2BD4: d <= 8'hC0; 15'h2BD5: d <= 8'hC0; 15'h2BD6: d <= 8'hC0; 15'h2BD7: d <= 8'hC0;
                15'h2BD8: d <= 8'hC0; 15'h2BD9: d <= 8'hC0; 15'h2BDA: d <= 8'hC0; 15'h2BDB: d <= 8'hC0;
                15'h2BDC: d <= 8'hC0; 15'h2BDD: d <= 8'hC0; 15'h2BDE: d <= 8'hC0; 15'h2BDF: d <= 8'hC0;
                15'h2BE0: d <= 8'hC0; 15'h2BE1: d <= 8'hC0; 15'h2BE2: d <= 8'hC0; 15'h2BE3: d <= 8'hC0;
                15'h2BE4: d <= 8'hC0; 15'h2BE5: d <= 8'hC0; 15'h2BE6: d <= 8'hC0; 15'h2BE7: d <= 8'hC0;
                15'h2BE8: d <= 8'hC0; 15'h2BE9: d <= 8'hC0; 15'h2BEA: d <= 8'hC0; 15'h2BEB: d <= 8'hC0;
                15'h2BEC: d <= 8'hC0; 15'h2BED: d <= 8'hC0; 15'h2BEE: d <= 8'hC0; 15'h2BEF: d <= 8'hC0;
                15'h2BF0: d <= 8'hC0; 15'h2BF1: d <= 8'hC0; 15'h2BF2: d <= 8'hC0; 15'h2BF3: d <= 8'hC0;
                15'h2BF4: d <= 8'hC0; 15'h2BF5: d <= 8'hC0; 15'h2BF6: d <= 8'hC0; 15'h2BF7: d <= 8'hC0;
                15'h2BF8: d <= 8'hC0; 15'h2BF9: d <= 8'hC0; 15'h2BFA: d <= 8'hC0; 15'h2BFB: d <= 8'hC0;
                15'h2BFC: d <= 8'hC0; 15'h2BFD: d <= 8'hC0; 15'h2BFE: d <= 8'hC0; 15'h2BFF: d <= 8'hC0;
                15'h2C00: d <= 8'hC0; 15'h2C01: d <= 8'hC0; 15'h2C02: d <= 8'hC0; 15'h2C03: d <= 8'hC0;
                15'h2C04: d <= 8'hC0; 15'h2C05: d <= 8'hC0; 15'h2C06: d <= 8'hC0; 15'h2C07: d <= 8'hC0;
                15'h2C08: d <= 8'hC0; 15'h2C09: d <= 8'hC0; 15'h2C0A: d <= 8'hC0; 15'h2C0B: d <= 8'hC0;
                15'h2C0C: d <= 8'hC0; 15'h2C0D: d <= 8'hC0; 15'h2C0E: d <= 8'hC0; 15'h2C0F: d <= 8'hC0;
                15'h2C10: d <= 8'hC0; 15'h2C11: d <= 8'hC0; 15'h2C12: d <= 8'hC0; 15'h2C13: d <= 8'hC0;
                15'h2C14: d <= 8'hC0; 15'h2C15: d <= 8'hC0; 15'h2C16: d <= 8'hC0; 15'h2C17: d <= 8'hC0;
                15'h2C18: d <= 8'hC0; 15'h2C19: d <= 8'hC0; 15'h2C1A: d <= 8'hC0; 15'h2C1B: d <= 8'hC0;
                15'h2C1C: d <= 8'hC0; 15'h2C1D: d <= 8'hC0; 15'h2C1E: d <= 8'hC0; 15'h2C1F: d <= 8'hC0;
                15'h2C20: d <= 8'hC0; 15'h2C21: d <= 8'hC0; 15'h2C22: d <= 8'hC0; 15'h2C23: d <= 8'hC0;
                15'h2C24: d <= 8'hC0; 15'h2C25: d <= 8'hC0; 15'h2C26: d <= 8'hC0; 15'h2C27: d <= 8'hC0;
                15'h2C28: d <= 8'hC0; 15'h2C29: d <= 8'hC0; 15'h2C2A: d <= 8'hC0; 15'h2C2B: d <= 8'hC0;
                15'h2C2C: d <= 8'hC0; 15'h2C2D: d <= 8'hC0; 15'h2C2E: d <= 8'hC0; 15'h2C2F: d <= 8'hC0;
                15'h2C30: d <= 8'hC0; 15'h2C31: d <= 8'hC0; 15'h2C32: d <= 8'hC0; 15'h2C33: d <= 8'hC0;
                15'h2C34: d <= 8'hC0; 15'h2C35: d <= 8'hC0; 15'h2C36: d <= 8'hC0; 15'h2C37: d <= 8'hC0;
                15'h2C38: d <= 8'hC0; 15'h2C39: d <= 8'hC0; 15'h2C3A: d <= 8'hC0; 15'h2C3B: d <= 8'hC0;
                15'h2C3C: d <= 8'hC0; 15'h2C3D: d <= 8'hC0; 15'h2C3E: d <= 8'hC0; 15'h2C3F: d <= 8'hC0;
                15'h2C40: d <= 8'hC0; 15'h2C41: d <= 8'hC0; 15'h2C42: d <= 8'hC0; 15'h2C43: d <= 8'hC0;
                15'h2C44: d <= 8'hC0; 15'h2C45: d <= 8'hC0; 15'h2C46: d <= 8'hC0; 15'h2C47: d <= 8'hC0;
                15'h2C48: d <= 8'hC0; 15'h2C49: d <= 8'hC0; 15'h2C4A: d <= 8'hC0; 15'h2C4B: d <= 8'hC0;
                15'h2C4C: d <= 8'hC0; 15'h2C4D: d <= 8'hC0; 15'h2C4E: d <= 8'hC0; 15'h2C4F: d <= 8'hC0;
                15'h2C50: d <= 8'hC0; 15'h2C51: d <= 8'hC0; 15'h2C52: d <= 8'hC0; 15'h2C53: d <= 8'hC0;
                15'h2C54: d <= 8'hC0; 15'h2C55: d <= 8'hC0; 15'h2C56: d <= 8'hC0; 15'h2C57: d <= 8'hC0;
                15'h2C58: d <= 8'hC0; 15'h2C59: d <= 8'hC0; 15'h2C5A: d <= 8'hC0; 15'h2C5B: d <= 8'hC0;
                15'h2C5C: d <= 8'hC0; 15'h2C5D: d <= 8'hC0; 15'h2C5E: d <= 8'hC0; 15'h2C5F: d <= 8'hC0;
                15'h2C60: d <= 8'hC0; 15'h2C61: d <= 8'hC0; 15'h2C62: d <= 8'hC0; 15'h2C63: d <= 8'hC0;
                15'h2C64: d <= 8'hC0; 15'h2C65: d <= 8'hC0; 15'h2C66: d <= 8'hC0; 15'h2C67: d <= 8'hC0;
                15'h2C68: d <= 8'hC0; 15'h2C69: d <= 8'hC0; 15'h2C6A: d <= 8'hC0; 15'h2C6B: d <= 8'hC0;
                15'h2C6C: d <= 8'hC0; 15'h2C6D: d <= 8'hC0; 15'h2C6E: d <= 8'hC0; 15'h2C6F: d <= 8'hC0;
                15'h2C70: d <= 8'hC0; 15'h2C71: d <= 8'hC0; 15'h2C72: d <= 8'hC0; 15'h2C73: d <= 8'hC0;
                15'h2C74: d <= 8'hC0; 15'h2C75: d <= 8'hC0; 15'h2C76: d <= 8'hC0; 15'h2C77: d <= 8'hC0;
                15'h2C78: d <= 8'hC0; 15'h2C79: d <= 8'hC0; 15'h2C7A: d <= 8'hC0; 15'h2C7B: d <= 8'hC0;
                15'h2C7C: d <= 8'hC0; 15'h2C7D: d <= 8'hC0; 15'h2C7E: d <= 8'hC0; 15'h2C7F: d <= 8'hC0;
                15'h2C80: d <= 8'hC0; 15'h2C81: d <= 8'hC0; 15'h2C82: d <= 8'hC0; 15'h2C83: d <= 8'hC0;
                15'h2C84: d <= 8'hC0; 15'h2C85: d <= 8'hC0; 15'h2C86: d <= 8'hC0; 15'h2C87: d <= 8'hC0;
                15'h2C88: d <= 8'hC0; 15'h2C89: d <= 8'hC0; 15'h2C8A: d <= 8'hC0; 15'h2C8B: d <= 8'hC0;
                15'h2C8C: d <= 8'hC0; 15'h2C8D: d <= 8'hC0; 15'h2C8E: d <= 8'hC0; 15'h2C8F: d <= 8'hC0;
                15'h2C90: d <= 8'hC0; 15'h2C91: d <= 8'hC0; 15'h2C92: d <= 8'hC0; 15'h2C93: d <= 8'hC0;
                15'h2C94: d <= 8'hC0; 15'h2C95: d <= 8'hC0; 15'h2C96: d <= 8'hC0; 15'h2C97: d <= 8'hC0;
                15'h2C98: d <= 8'hC0; 15'h2C99: d <= 8'hC0; 15'h2C9A: d <= 8'hC0; 15'h2C9B: d <= 8'hC0;
                15'h2C9C: d <= 8'hC0; 15'h2C9D: d <= 8'hC0; 15'h2C9E: d <= 8'hC0; 15'h2C9F: d <= 8'hC0;
                15'h2CA0: d <= 8'hC0; 15'h2CA1: d <= 8'hC0; 15'h2CA2: d <= 8'hC0; 15'h2CA3: d <= 8'hC0;
                15'h2CA4: d <= 8'hC0; 15'h2CA5: d <= 8'hC0; 15'h2CA6: d <= 8'hC0; 15'h2CA7: d <= 8'hC0;
                15'h2CA8: d <= 8'hC0; 15'h2CA9: d <= 8'hC0; 15'h2CAA: d <= 8'hC0; 15'h2CAB: d <= 8'hC0;
                15'h2CAC: d <= 8'hC0; 15'h2CAD: d <= 8'hC0; 15'h2CAE: d <= 8'hC0; 15'h2CAF: d <= 8'hC0;
                15'h2CB0: d <= 8'hC0; 15'h2CB1: d <= 8'hC0; 15'h2CB2: d <= 8'hC0; 15'h2CB3: d <= 8'hC0;
                15'h2CB4: d <= 8'hC0; 15'h2CB5: d <= 8'hC0; 15'h2CB6: d <= 8'hC0; 15'h2CB7: d <= 8'hC0;
                15'h2CB8: d <= 8'hC0; 15'h2CB9: d <= 8'hC0; 15'h2CBA: d <= 8'hC0; 15'h2CBB: d <= 8'hC0;
                15'h2CBC: d <= 8'hC0; 15'h2CBD: d <= 8'hC0; 15'h2CBE: d <= 8'hC0; 15'h2CBF: d <= 8'hC0;
                15'h2CC0: d <= 8'hC0; 15'h2CC1: d <= 8'hC0; 15'h2CC2: d <= 8'hC0; 15'h2CC3: d <= 8'hC0;
                15'h2CC4: d <= 8'hC0; 15'h2CC5: d <= 8'hC0; 15'h2CC6: d <= 8'hC0; 15'h2CC7: d <= 8'hC0;
                15'h2CC8: d <= 8'hC0; 15'h2CC9: d <= 8'hC0; 15'h2CCA: d <= 8'hC0; 15'h2CCB: d <= 8'hC0;
                15'h2CCC: d <= 8'hC0; 15'h2CCD: d <= 8'hC0; 15'h2CCE: d <= 8'hC0; 15'h2CCF: d <= 8'hC0;
                15'h2CD0: d <= 8'hC0; 15'h2CD1: d <= 8'hC0; 15'h2CD2: d <= 8'hC0; 15'h2CD3: d <= 8'hC0;
                15'h2CD4: d <= 8'hC0; 15'h2CD5: d <= 8'hC0; 15'h2CD6: d <= 8'hC0; 15'h2CD7: d <= 8'hC0;
                15'h2CD8: d <= 8'hC0; 15'h2CD9: d <= 8'hC0; 15'h2CDA: d <= 8'hC0; 15'h2CDB: d <= 8'hC0;
                15'h2CDC: d <= 8'hC0; 15'h2CDD: d <= 8'hC0; 15'h2CDE: d <= 8'hC0; 15'h2CDF: d <= 8'hC0;
                15'h2CE0: d <= 8'hC0; 15'h2CE1: d <= 8'hC0; 15'h2CE2: d <= 8'hC0; 15'h2CE3: d <= 8'hC0;
                15'h2CE4: d <= 8'hC0; 15'h2CE5: d <= 8'hC0; 15'h2CE6: d <= 8'hC0; 15'h2CE7: d <= 8'hC0;
                15'h2CE8: d <= 8'hC0; 15'h2CE9: d <= 8'hC0; 15'h2CEA: d <= 8'hC0; 15'h2CEB: d <= 8'hC0;
                15'h2CEC: d <= 8'hC0; 15'h2CED: d <= 8'hC0; 15'h2CEE: d <= 8'hC0; 15'h2CEF: d <= 8'hC0;
                15'h2CF0: d <= 8'hC0; 15'h2CF1: d <= 8'hC0; 15'h2CF2: d <= 8'hC0; 15'h2CF3: d <= 8'hC0;
                15'h2CF4: d <= 8'hC0; 15'h2CF5: d <= 8'hC0; 15'h2CF6: d <= 8'hC0; 15'h2CF7: d <= 8'hC0;
                15'h2CF8: d <= 8'hC0; 15'h2CF9: d <= 8'hC0; 15'h2CFA: d <= 8'hC0; 15'h2CFB: d <= 8'hC0;
                15'h2CFC: d <= 8'hC0; 15'h2CFD: d <= 8'hC0; 15'h2CFE: d <= 8'hC0; 15'h2CFF: d <= 8'hC0;
                15'h2D00: d <= 8'hC0; 15'h2D01: d <= 8'hC0; 15'h2D02: d <= 8'hC0; 15'h2D03: d <= 8'hC0;
                15'h2D04: d <= 8'hC0; 15'h2D05: d <= 8'hC0; 15'h2D06: d <= 8'hC0; 15'h2D07: d <= 8'hC0;
                15'h2D08: d <= 8'hC0; 15'h2D09: d <= 8'hC0; 15'h2D0A: d <= 8'hC0; 15'h2D0B: d <= 8'hC0;
                15'h2D0C: d <= 8'hC0; 15'h2D0D: d <= 8'hC0; 15'h2D0E: d <= 8'hC0; 15'h2D0F: d <= 8'hC0;
                15'h2D10: d <= 8'hC0; 15'h2D11: d <= 8'hC0; 15'h2D12: d <= 8'hC0; 15'h2D13: d <= 8'hC0;
                15'h2D14: d <= 8'hC0; 15'h2D15: d <= 8'hC0; 15'h2D16: d <= 8'hC0; 15'h2D17: d <= 8'hC0;
                15'h2D18: d <= 8'hC0; 15'h2D19: d <= 8'hC0; 15'h2D1A: d <= 8'hC0; 15'h2D1B: d <= 8'hC0;
                15'h2D1C: d <= 8'hC0; 15'h2D1D: d <= 8'hC0; 15'h2D1E: d <= 8'hC0; 15'h2D1F: d <= 8'hC0;
                15'h2D20: d <= 8'hC0; 15'h2D21: d <= 8'hC0; 15'h2D22: d <= 8'hC0; 15'h2D23: d <= 8'hC0;
                15'h2D24: d <= 8'hC0; 15'h2D25: d <= 8'hC0; 15'h2D26: d <= 8'hC0; 15'h2D27: d <= 8'hC0;
                15'h2D28: d <= 8'hC0; 15'h2D29: d <= 8'hC0; 15'h2D2A: d <= 8'hC0; 15'h2D2B: d <= 8'hC0;
                15'h2D2C: d <= 8'hC0; 15'h2D2D: d <= 8'hC0; 15'h2D2E: d <= 8'hC0; 15'h2D2F: d <= 8'hC0;
                15'h2D30: d <= 8'hC0; 15'h2D31: d <= 8'hC0; 15'h2D32: d <= 8'hC0; 15'h2D33: d <= 8'hC0;
                15'h2D34: d <= 8'hC0; 15'h2D35: d <= 8'hC0; 15'h2D36: d <= 8'hC0; 15'h2D37: d <= 8'hC0;
                15'h2D38: d <= 8'hC0; 15'h2D39: d <= 8'hC0; 15'h2D3A: d <= 8'hC0; 15'h2D3B: d <= 8'hC0;
                15'h2D3C: d <= 8'hC0; 15'h2D3D: d <= 8'hC0; 15'h2D3E: d <= 8'hC0; 15'h2D3F: d <= 8'hC0;
                15'h2D40: d <= 8'hC0; 15'h2D41: d <= 8'hC0; 15'h2D42: d <= 8'hC0; 15'h2D43: d <= 8'hC0;
                15'h2D44: d <= 8'hC0; 15'h2D45: d <= 8'hC0; 15'h2D46: d <= 8'hC0; 15'h2D47: d <= 8'hC0;
                15'h2D48: d <= 8'hC0; 15'h2D49: d <= 8'hC0; 15'h2D4A: d <= 8'hC0; 15'h2D4B: d <= 8'hC0;
                15'h2D4C: d <= 8'hC0; 15'h2D4D: d <= 8'hC0; 15'h2D4E: d <= 8'hC0; 15'h2D4F: d <= 8'hC0;
                15'h2D50: d <= 8'hC0; 15'h2D51: d <= 8'hC0; 15'h2D52: d <= 8'hC0; 15'h2D53: d <= 8'hC0;
                15'h2D54: d <= 8'hC0; 15'h2D55: d <= 8'hC0; 15'h2D56: d <= 8'hC0; 15'h2D57: d <= 8'hC0;
                15'h2D58: d <= 8'hC0; 15'h2D59: d <= 8'hC0; 15'h2D5A: d <= 8'hC0; 15'h2D5B: d <= 8'hC0;
                15'h2D5C: d <= 8'hC0; 15'h2D5D: d <= 8'hC0; 15'h2D5E: d <= 8'hC0; 15'h2D5F: d <= 8'hC0;
                15'h2D60: d <= 8'hC0; 15'h2D61: d <= 8'hC0; 15'h2D62: d <= 8'hC0; 15'h2D63: d <= 8'hC0;
                15'h2D64: d <= 8'hC0; 15'h2D65: d <= 8'hC0; 15'h2D66: d <= 8'hC0; 15'h2D67: d <= 8'hC0;
                15'h2D68: d <= 8'hC0; 15'h2D69: d <= 8'hC0; 15'h2D6A: d <= 8'hC0; 15'h2D6B: d <= 8'hC0;
                15'h2D6C: d <= 8'hC0; 15'h2D6D: d <= 8'hC0; 15'h2D6E: d <= 8'hC0; 15'h2D6F: d <= 8'hC0;
                15'h2D70: d <= 8'hC0; 15'h2D71: d <= 8'hC0; 15'h2D72: d <= 8'hC0; 15'h2D73: d <= 8'hC0;
                15'h2D74: d <= 8'hC0; 15'h2D75: d <= 8'hC0; 15'h2D76: d <= 8'hC0; 15'h2D77: d <= 8'hC0;
                15'h2D78: d <= 8'hC0; 15'h2D79: d <= 8'hC0; 15'h2D7A: d <= 8'hC0; 15'h2D7B: d <= 8'hC0;
                15'h2D7C: d <= 8'hC0; 15'h2D7D: d <= 8'hC0; 15'h2D7E: d <= 8'hC0; 15'h2D7F: d <= 8'hC0;
                15'h2D80: d <= 8'hC0; 15'h2D81: d <= 8'hC0; 15'h2D82: d <= 8'hC0; 15'h2D83: d <= 8'hC0;
                15'h2D84: d <= 8'hC0; 15'h2D85: d <= 8'hC0; 15'h2D86: d <= 8'hC0; 15'h2D87: d <= 8'hC0;
                15'h2D88: d <= 8'hC0; 15'h2D89: d <= 8'hC0; 15'h2D8A: d <= 8'hC0; 15'h2D8B: d <= 8'hC0;
                15'h2D8C: d <= 8'hC0; 15'h2D8D: d <= 8'hC0; 15'h2D8E: d <= 8'hC0; 15'h2D8F: d <= 8'hC0;
                15'h2D90: d <= 8'hC0; 15'h2D91: d <= 8'hC0; 15'h2D92: d <= 8'hC0; 15'h2D93: d <= 8'hC0;
                15'h2D94: d <= 8'hC0; 15'h2D95: d <= 8'hC0; 15'h2D96: d <= 8'hC0; 15'h2D97: d <= 8'hC0;
                15'h2D98: d <= 8'hC0; 15'h2D99: d <= 8'hC0; 15'h2D9A: d <= 8'hC0; 15'h2D9B: d <= 8'hC0;
                15'h2D9C: d <= 8'hC0; 15'h2D9D: d <= 8'hC0; 15'h2D9E: d <= 8'hC0; 15'h2D9F: d <= 8'hC0;
                15'h2DA0: d <= 8'hC0; 15'h2DA1: d <= 8'hC0; 15'h2DA2: d <= 8'hC0; 15'h2DA3: d <= 8'hC0;
                15'h2DA4: d <= 8'hC0; 15'h2DA5: d <= 8'hC0; 15'h2DA6: d <= 8'hC0; 15'h2DA7: d <= 8'hC0;
                15'h2DA8: d <= 8'hC0; 15'h2DA9: d <= 8'hC0; 15'h2DAA: d <= 8'hC0; 15'h2DAB: d <= 8'hC0;
                15'h2DAC: d <= 8'hC0; 15'h2DAD: d <= 8'hC0; 15'h2DAE: d <= 8'hC0; 15'h2DAF: d <= 8'hC0;
                15'h2DB0: d <= 8'hC0; 15'h2DB1: d <= 8'hC0; 15'h2DB2: d <= 8'hC0; 15'h2DB3: d <= 8'hC0;
                15'h2DB4: d <= 8'hC0; 15'h2DB5: d <= 8'hC0; 15'h2DB6: d <= 8'hC0; 15'h2DB7: d <= 8'hC0;
                15'h2DB8: d <= 8'hC0; 15'h2DB9: d <= 8'hC0; 15'h2DBA: d <= 8'hC0; 15'h2DBB: d <= 8'hC0;
                15'h2DBC: d <= 8'hC0; 15'h2DBD: d <= 8'hC0; 15'h2DBE: d <= 8'hC0; 15'h2DBF: d <= 8'hC0;
                15'h2DC0: d <= 8'hC0; 15'h2DC1: d <= 8'hC0; 15'h2DC2: d <= 8'hC0; 15'h2DC3: d <= 8'hC0;
                15'h2DC4: d <= 8'hC0; 15'h2DC5: d <= 8'hC0; 15'h2DC6: d <= 8'hC0; 15'h2DC7: d <= 8'hC0;
                15'h2DC8: d <= 8'hC0; 15'h2DC9: d <= 8'hC0; 15'h2DCA: d <= 8'hC0; 15'h2DCB: d <= 8'hC0;
                15'h2DCC: d <= 8'hC0; 15'h2DCD: d <= 8'hC0; 15'h2DCE: d <= 8'hC0; 15'h2DCF: d <= 8'hC0;
                15'h2DD0: d <= 8'hC0; 15'h2DD1: d <= 8'hC0; 15'h2DD2: d <= 8'hC0; 15'h2DD3: d <= 8'hC0;
                15'h2DD4: d <= 8'hC0; 15'h2DD5: d <= 8'hC0; 15'h2DD6: d <= 8'hC0; 15'h2DD7: d <= 8'hC0;
                15'h2DD8: d <= 8'hC0; 15'h2DD9: d <= 8'hC0; 15'h2DDA: d <= 8'hC0; 15'h2DDB: d <= 8'hC0;
                15'h2DDC: d <= 8'hC0; 15'h2DDD: d <= 8'hC0; 15'h2DDE: d <= 8'hC0; 15'h2DDF: d <= 8'hC0;
                15'h2DE0: d <= 8'hC0; 15'h2DE1: d <= 8'hC0; 15'h2DE2: d <= 8'hC0; 15'h2DE3: d <= 8'hC0;
                15'h2DE4: d <= 8'hC0; 15'h2DE5: d <= 8'hC0; 15'h2DE6: d <= 8'hC0; 15'h2DE7: d <= 8'hC0;
                15'h2DE8: d <= 8'hC0; 15'h2DE9: d <= 8'hC0; 15'h2DEA: d <= 8'hC0; 15'h2DEB: d <= 8'hC0;
                15'h2DEC: d <= 8'hC0; 15'h2DED: d <= 8'hC0; 15'h2DEE: d <= 8'hC0; 15'h2DEF: d <= 8'hC0;
                15'h2DF0: d <= 8'hC0; 15'h2DF1: d <= 8'hC0; 15'h2DF2: d <= 8'hC0; 15'h2DF3: d <= 8'hC0;
                15'h2DF4: d <= 8'hC0; 15'h2DF5: d <= 8'hC0; 15'h2DF6: d <= 8'hC0; 15'h2DF7: d <= 8'hC0;
                15'h2DF8: d <= 8'hC0; 15'h2DF9: d <= 8'hC0; 15'h2DFA: d <= 8'hC0; 15'h2DFB: d <= 8'hC0;
                15'h2DFC: d <= 8'hC0; 15'h2DFD: d <= 8'hC0; 15'h2DFE: d <= 8'hC0; 15'h2DFF: d <= 8'hC0;
                15'h2E00: d <= 8'hC0; 15'h2E01: d <= 8'hC0; 15'h2E02: d <= 8'hC0; 15'h2E03: d <= 8'hC0;
                15'h2E04: d <= 8'hC0; 15'h2E05: d <= 8'hC0; 15'h2E06: d <= 8'hC0; 15'h2E07: d <= 8'hC0;
                15'h2E08: d <= 8'hC0; 15'h2E09: d <= 8'hC0; 15'h2E0A: d <= 8'hC0; 15'h2E0B: d <= 8'hC0;
                15'h2E0C: d <= 8'hC0; 15'h2E0D: d <= 8'hC0; 15'h2E0E: d <= 8'hC0; 15'h2E0F: d <= 8'hC0;
                15'h2E10: d <= 8'hC0; 15'h2E11: d <= 8'hC0; 15'h2E12: d <= 8'hC0; 15'h2E13: d <= 8'hC0;
                15'h2E14: d <= 8'hC0; 15'h2E15: d <= 8'hC0; 15'h2E16: d <= 8'hC0; 15'h2E17: d <= 8'hC0;
                15'h2E18: d <= 8'hC0; 15'h2E19: d <= 8'hC0; 15'h2E1A: d <= 8'hC0; 15'h2E1B: d <= 8'hC0;
                15'h2E1C: d <= 8'hC0; 15'h2E1D: d <= 8'hC0; 15'h2E1E: d <= 8'hC0; 15'h2E1F: d <= 8'hC0;
                15'h2E20: d <= 8'hC0; 15'h2E21: d <= 8'hC0; 15'h2E22: d <= 8'hC0; 15'h2E23: d <= 8'hC0;
                15'h2E24: d <= 8'hC0; 15'h2E25: d <= 8'hC0; 15'h2E26: d <= 8'hC0; 15'h2E27: d <= 8'hC0;
                15'h2E28: d <= 8'hC0; 15'h2E29: d <= 8'hC0; 15'h2E2A: d <= 8'hC0; 15'h2E2B: d <= 8'hC0;
                15'h2E2C: d <= 8'hC0; 15'h2E2D: d <= 8'hC0; 15'h2E2E: d <= 8'hC0; 15'h2E2F: d <= 8'hC0;
                15'h2E30: d <= 8'hC0; 15'h2E31: d <= 8'hC0; 15'h2E32: d <= 8'hC0; 15'h2E33: d <= 8'hC0;
                15'h2E34: d <= 8'hC0; 15'h2E35: d <= 8'hC0; 15'h2E36: d <= 8'hC0; 15'h2E37: d <= 8'hC0;
                15'h2E38: d <= 8'hC0; 15'h2E39: d <= 8'hC0; 15'h2E3A: d <= 8'hC0; 15'h2E3B: d <= 8'hC0;
                15'h2E3C: d <= 8'hC0; 15'h2E3D: d <= 8'hC0; 15'h2E3E: d <= 8'hC0; 15'h2E3F: d <= 8'hC0;
                15'h2E40: d <= 8'hC0; 15'h2E41: d <= 8'hC0; 15'h2E42: d <= 8'hC0; 15'h2E43: d <= 8'hC0;
                15'h2E44: d <= 8'hC0; 15'h2E45: d <= 8'hC0; 15'h2E46: d <= 8'hC0; 15'h2E47: d <= 8'hC0;
                15'h2E48: d <= 8'hC0; 15'h2E49: d <= 8'hC0; 15'h2E4A: d <= 8'hC0; 15'h2E4B: d <= 8'hC0;
                15'h2E4C: d <= 8'hC0; 15'h2E4D: d <= 8'hC0; 15'h2E4E: d <= 8'hC0; 15'h2E4F: d <= 8'hC0;
                15'h2E50: d <= 8'hC0; 15'h2E51: d <= 8'hC0; 15'h2E52: d <= 8'hC0; 15'h2E53: d <= 8'hC0;
                15'h2E54: d <= 8'hC0; 15'h2E55: d <= 8'hC0; 15'h2E56: d <= 8'hC0; 15'h2E57: d <= 8'hC0;
                15'h2E58: d <= 8'hC0; 15'h2E59: d <= 8'hC0; 15'h2E5A: d <= 8'hC0; 15'h2E5B: d <= 8'hC0;
                15'h2E5C: d <= 8'hC0; 15'h2E5D: d <= 8'hC0; 15'h2E5E: d <= 8'hC0; 15'h2E5F: d <= 8'hC0;
                15'h2E60: d <= 8'hC0; 15'h2E61: d <= 8'hC0; 15'h2E62: d <= 8'hC0; 15'h2E63: d <= 8'hC0;
                15'h2E64: d <= 8'hC0; 15'h2E65: d <= 8'hC0; 15'h2E66: d <= 8'hC0; 15'h2E67: d <= 8'hC0;
                15'h2E68: d <= 8'hC0; 15'h2E69: d <= 8'hC0; 15'h2E6A: d <= 8'hC0; 15'h2E6B: d <= 8'hC0;
                15'h2E6C: d <= 8'hC0; 15'h2E6D: d <= 8'hC0; 15'h2E6E: d <= 8'hC0; 15'h2E6F: d <= 8'hC0;
                15'h2E70: d <= 8'hC0; 15'h2E71: d <= 8'hC0; 15'h2E72: d <= 8'hC0; 15'h2E73: d <= 8'hC0;
                15'h2E74: d <= 8'hC0; 15'h2E75: d <= 8'hC0; 15'h2E76: d <= 8'hC0; 15'h2E77: d <= 8'hC0;
                15'h2E78: d <= 8'hC0; 15'h2E79: d <= 8'hC0; 15'h2E7A: d <= 8'hC0; 15'h2E7B: d <= 8'hC0;
                15'h2E7C: d <= 8'hC0; 15'h2E7D: d <= 8'hC0; 15'h2E7E: d <= 8'hC0; 15'h2E7F: d <= 8'hC0;
                15'h2E80: d <= 8'hC0; 15'h2E81: d <= 8'hC0; 15'h2E82: d <= 8'hC0; 15'h2E83: d <= 8'hC0;
                15'h2E84: d <= 8'hC0; 15'h2E85: d <= 8'hC0; 15'h2E86: d <= 8'hC0; 15'h2E87: d <= 8'hC0;
                15'h2E88: d <= 8'hC0; 15'h2E89: d <= 8'hC0; 15'h2E8A: d <= 8'hC0; 15'h2E8B: d <= 8'hC0;
                15'h2E8C: d <= 8'hC0; 15'h2E8D: d <= 8'hC0; 15'h2E8E: d <= 8'hC0; 15'h2E8F: d <= 8'hC0;
                15'h2E90: d <= 8'hC0; 15'h2E91: d <= 8'hC0; 15'h2E92: d <= 8'hC0; 15'h2E93: d <= 8'hC0;
                15'h2E94: d <= 8'hC0; 15'h2E95: d <= 8'hC0; 15'h2E96: d <= 8'hC0; 15'h2E97: d <= 8'hC0;
                15'h2E98: d <= 8'hC0; 15'h2E99: d <= 8'hC0; 15'h2E9A: d <= 8'hC0; 15'h2E9B: d <= 8'hC0;
                15'h2E9C: d <= 8'hC0; 15'h2E9D: d <= 8'hC0; 15'h2E9E: d <= 8'hC0; 15'h2E9F: d <= 8'hC0;
                15'h2EA0: d <= 8'hC0; 15'h2EA1: d <= 8'hC0; 15'h2EA2: d <= 8'hC0; 15'h2EA3: d <= 8'hC0;
                15'h2EA4: d <= 8'hC0; 15'h2EA5: d <= 8'hC0; 15'h2EA6: d <= 8'hC0; 15'h2EA7: d <= 8'hC0;
                15'h2EA8: d <= 8'hC0; 15'h2EA9: d <= 8'hC0; 15'h2EAA: d <= 8'hC0; 15'h2EAB: d <= 8'hC0;
                15'h2EAC: d <= 8'hC0; 15'h2EAD: d <= 8'hC0; 15'h2EAE: d <= 8'hC0; 15'h2EAF: d <= 8'hC0;
                15'h2EB0: d <= 8'hC0; 15'h2EB1: d <= 8'hC0; 15'h2EB2: d <= 8'hC0; 15'h2EB3: d <= 8'hC0;
                15'h2EB4: d <= 8'hC0; 15'h2EB5: d <= 8'hC0; 15'h2EB6: d <= 8'hC0; 15'h2EB7: d <= 8'hC0;
                15'h2EB8: d <= 8'hC0; 15'h2EB9: d <= 8'hC0; 15'h2EBA: d <= 8'hC0; 15'h2EBB: d <= 8'hC0;
                15'h2EBC: d <= 8'hC0; 15'h2EBD: d <= 8'hC0; 15'h2EBE: d <= 8'hC0; 15'h2EBF: d <= 8'hC0;
                15'h2EC0: d <= 8'hC0; 15'h2EC1: d <= 8'hC0; 15'h2EC2: d <= 8'hC0; 15'h2EC3: d <= 8'hC0;
                15'h2EC4: d <= 8'hC0; 15'h2EC5: d <= 8'hC0; 15'h2EC6: d <= 8'hC0; 15'h2EC7: d <= 8'hC0;
                15'h2EC8: d <= 8'hC0; 15'h2EC9: d <= 8'hC0; 15'h2ECA: d <= 8'hC0; 15'h2ECB: d <= 8'hC0;
                15'h2ECC: d <= 8'hC0; 15'h2ECD: d <= 8'hC0; 15'h2ECE: d <= 8'hC0; 15'h2ECF: d <= 8'hC0;
                15'h2ED0: d <= 8'hC0; 15'h2ED1: d <= 8'hC0; 15'h2ED2: d <= 8'hC0; 15'h2ED3: d <= 8'hC0;
                15'h2ED4: d <= 8'hC0; 15'h2ED5: d <= 8'hC0; 15'h2ED6: d <= 8'hC0; 15'h2ED7: d <= 8'hC0;
                15'h2ED8: d <= 8'hC0; 15'h2ED9: d <= 8'hC0; 15'h2EDA: d <= 8'hC0; 15'h2EDB: d <= 8'hC0;
                15'h2EDC: d <= 8'hC0; 15'h2EDD: d <= 8'hC0; 15'h2EDE: d <= 8'hC0; 15'h2EDF: d <= 8'hC0;
                15'h2EE0: d <= 8'hC0; 15'h2EE1: d <= 8'hC0; 15'h2EE2: d <= 8'hC0; 15'h2EE3: d <= 8'hC0;
                15'h2EE4: d <= 8'hC0; 15'h2EE5: d <= 8'hC0; 15'h2EE6: d <= 8'hC0; 15'h2EE7: d <= 8'hC0;
                15'h2EE8: d <= 8'hC0; 15'h2EE9: d <= 8'hC0; 15'h2EEA: d <= 8'hC0; 15'h2EEB: d <= 8'hC0;
                15'h2EEC: d <= 8'hC0; 15'h2EED: d <= 8'hC0; 15'h2EEE: d <= 8'hC0; 15'h2EEF: d <= 8'hC0;
                15'h2EF0: d <= 8'hC0; 15'h2EF1: d <= 8'hC0; 15'h2EF2: d <= 8'hC0; 15'h2EF3: d <= 8'hC0;
                15'h2EF4: d <= 8'hC0; 15'h2EF5: d <= 8'hC0; 15'h2EF6: d <= 8'hC0; 15'h2EF7: d <= 8'hC0;
                15'h2EF8: d <= 8'hC0; 15'h2EF9: d <= 8'hC0; 15'h2EFA: d <= 8'hC0; 15'h2EFB: d <= 8'hC0;
                15'h2EFC: d <= 8'hC0; 15'h2EFD: d <= 8'hC0; 15'h2EFE: d <= 8'hC0; 15'h2EFF: d <= 8'hC0;
                15'h2F00: d <= 8'hC0; 15'h2F01: d <= 8'hC0; 15'h2F02: d <= 8'hC0; 15'h2F03: d <= 8'hC0;
                15'h2F04: d <= 8'hC0; 15'h2F05: d <= 8'hC0; 15'h2F06: d <= 8'hC0; 15'h2F07: d <= 8'hC0;
                15'h2F08: d <= 8'hC0; 15'h2F09: d <= 8'hC0; 15'h2F0A: d <= 8'hC0; 15'h2F0B: d <= 8'hC0;
                15'h2F0C: d <= 8'hC0; 15'h2F0D: d <= 8'hC0; 15'h2F0E: d <= 8'hC0; 15'h2F0F: d <= 8'hC0;
                15'h2F10: d <= 8'hC0; 15'h2F11: d <= 8'hC0; 15'h2F12: d <= 8'hC0; 15'h2F13: d <= 8'hC0;
                15'h2F14: d <= 8'hC0; 15'h2F15: d <= 8'hC0; 15'h2F16: d <= 8'hC0; 15'h2F17: d <= 8'hC0;
                15'h2F18: d <= 8'hC0; 15'h2F19: d <= 8'hC0; 15'h2F1A: d <= 8'hC0; 15'h2F1B: d <= 8'hC0;
                15'h2F1C: d <= 8'hC0; 15'h2F1D: d <= 8'hC0; 15'h2F1E: d <= 8'hC0; 15'h2F1F: d <= 8'hC0;
                15'h2F20: d <= 8'hC0; 15'h2F21: d <= 8'hC0; 15'h2F22: d <= 8'hC0; 15'h2F23: d <= 8'hC0;
                15'h2F24: d <= 8'hC0; 15'h2F25: d <= 8'hC0; 15'h2F26: d <= 8'hC0; 15'h2F27: d <= 8'hC0;
                15'h2F28: d <= 8'hC0; 15'h2F29: d <= 8'hC0; 15'h2F2A: d <= 8'hC0; 15'h2F2B: d <= 8'hC0;
                15'h2F2C: d <= 8'hC0; 15'h2F2D: d <= 8'hC0; 15'h2F2E: d <= 8'hC0; 15'h2F2F: d <= 8'hC0;
                15'h2F30: d <= 8'hC0; 15'h2F31: d <= 8'hC0; 15'h2F32: d <= 8'hC0; 15'h2F33: d <= 8'hC0;
                15'h2F34: d <= 8'hC0; 15'h2F35: d <= 8'hC0; 15'h2F36: d <= 8'hC0; 15'h2F37: d <= 8'hC0;
                15'h2F38: d <= 8'hC0; 15'h2F39: d <= 8'hC0; 15'h2F3A: d <= 8'hC0; 15'h2F3B: d <= 8'hC0;
                15'h2F3C: d <= 8'hC0; 15'h2F3D: d <= 8'hC0; 15'h2F3E: d <= 8'hC0; 15'h2F3F: d <= 8'hC0;
                15'h2F40: d <= 8'hC0; 15'h2F41: d <= 8'hC0; 15'h2F42: d <= 8'hC0; 15'h2F43: d <= 8'hC0;
                15'h2F44: d <= 8'hC0; 15'h2F45: d <= 8'hC0; 15'h2F46: d <= 8'hC0; 15'h2F47: d <= 8'hC0;
                15'h2F48: d <= 8'hC0; 15'h2F49: d <= 8'hC0; 15'h2F4A: d <= 8'hC0; 15'h2F4B: d <= 8'hC0;
                15'h2F4C: d <= 8'hC0; 15'h2F4D: d <= 8'hC0; 15'h2F4E: d <= 8'hC0; 15'h2F4F: d <= 8'hC0;
                15'h2F50: d <= 8'hC0; 15'h2F51: d <= 8'hC0; 15'h2F52: d <= 8'hC0; 15'h2F53: d <= 8'hC0;
                15'h2F54: d <= 8'hC0; 15'h2F55: d <= 8'hC0; 15'h2F56: d <= 8'hC0; 15'h2F57: d <= 8'hC0;
                15'h2F58: d <= 8'hC0; 15'h2F59: d <= 8'hC0; 15'h2F5A: d <= 8'hC0; 15'h2F5B: d <= 8'hC0;
                15'h2F5C: d <= 8'hC0; 15'h2F5D: d <= 8'hC0; 15'h2F5E: d <= 8'hC0; 15'h2F5F: d <= 8'hC0;
                15'h2F60: d <= 8'hC0; 15'h2F61: d <= 8'hC0; 15'h2F62: d <= 8'hC0; 15'h2F63: d <= 8'hC0;
                15'h2F64: d <= 8'hC0; 15'h2F65: d <= 8'hC0; 15'h2F66: d <= 8'hC0; 15'h2F67: d <= 8'hC0;
                15'h2F68: d <= 8'hC0; 15'h2F69: d <= 8'hC0; 15'h2F6A: d <= 8'hC0; 15'h2F6B: d <= 8'hC0;
                15'h2F6C: d <= 8'hC0; 15'h2F6D: d <= 8'hC0; 15'h2F6E: d <= 8'hC0; 15'h2F6F: d <= 8'hC0;
                15'h2F70: d <= 8'hC0; 15'h2F71: d <= 8'hC0; 15'h2F72: d <= 8'hC0; 15'h2F73: d <= 8'hC0;
                15'h2F74: d <= 8'hC0; 15'h2F75: d <= 8'hC0; 15'h2F76: d <= 8'hC0; 15'h2F77: d <= 8'hC0;
                15'h2F78: d <= 8'hC0; 15'h2F79: d <= 8'hC0; 15'h2F7A: d <= 8'hC0; 15'h2F7B: d <= 8'hC0;
                15'h2F7C: d <= 8'hC0; 15'h2F7D: d <= 8'hC0; 15'h2F7E: d <= 8'hC0; 15'h2F7F: d <= 8'hC0;
                15'h2F80: d <= 8'hC0; 15'h2F81: d <= 8'hC0; 15'h2F82: d <= 8'hC0; 15'h2F83: d <= 8'hC0;
                15'h2F84: d <= 8'hC0; 15'h2F85: d <= 8'hC0; 15'h2F86: d <= 8'hC0; 15'h2F87: d <= 8'hC0;
                15'h2F88: d <= 8'hC0; 15'h2F89: d <= 8'hC0; 15'h2F8A: d <= 8'hC0; 15'h2F8B: d <= 8'hC0;
                15'h2F8C: d <= 8'hC0; 15'h2F8D: d <= 8'hC0; 15'h2F8E: d <= 8'hC0; 15'h2F8F: d <= 8'hC0;
                15'h2F90: d <= 8'hC0; 15'h2F91: d <= 8'hC0; 15'h2F92: d <= 8'hC0; 15'h2F93: d <= 8'hC0;
                15'h2F94: d <= 8'hC0; 15'h2F95: d <= 8'hC0; 15'h2F96: d <= 8'hC0; 15'h2F97: d <= 8'hC0;
                15'h2F98: d <= 8'hC0; 15'h2F99: d <= 8'hC0; 15'h2F9A: d <= 8'hC0; 15'h2F9B: d <= 8'hC0;
                15'h2F9C: d <= 8'hC0; 15'h2F9D: d <= 8'hC0; 15'h2F9E: d <= 8'hC0; 15'h2F9F: d <= 8'hC0;
                15'h2FA0: d <= 8'hC0; 15'h2FA1: d <= 8'hC0; 15'h2FA2: d <= 8'hC0; 15'h2FA3: d <= 8'hC0;
                15'h2FA4: d <= 8'hC0; 15'h2FA5: d <= 8'hC0; 15'h2FA6: d <= 8'hC0; 15'h2FA7: d <= 8'hC0;
                15'h2FA8: d <= 8'hC0; 15'h2FA9: d <= 8'hC0; 15'h2FAA: d <= 8'hC0; 15'h2FAB: d <= 8'hC0;
                15'h2FAC: d <= 8'hC0; 15'h2FAD: d <= 8'hC0; 15'h2FAE: d <= 8'hC0; 15'h2FAF: d <= 8'hC0;
                15'h2FB0: d <= 8'hC0; 15'h2FB1: d <= 8'hC0; 15'h2FB2: d <= 8'hC0; 15'h2FB3: d <= 8'hC0;
                15'h2FB4: d <= 8'hC0; 15'h2FB5: d <= 8'hC0; 15'h2FB6: d <= 8'hC0; 15'h2FB7: d <= 8'hC0;
                15'h2FB8: d <= 8'hC0; 15'h2FB9: d <= 8'hC0; 15'h2FBA: d <= 8'hC0; 15'h2FBB: d <= 8'hC0;
                15'h2FBC: d <= 8'hC0; 15'h2FBD: d <= 8'hC0; 15'h2FBE: d <= 8'hC0; 15'h2FBF: d <= 8'hC0;
                15'h2FC0: d <= 8'hC0; 15'h2FC1: d <= 8'hC0; 15'h2FC2: d <= 8'hC0; 15'h2FC3: d <= 8'hC0;
                15'h2FC4: d <= 8'hC0; 15'h2FC5: d <= 8'hC0; 15'h2FC6: d <= 8'hC0; 15'h2FC7: d <= 8'hC0;
                15'h2FC8: d <= 8'hC0; 15'h2FC9: d <= 8'hC0; 15'h2FCA: d <= 8'hC0; 15'h2FCB: d <= 8'hC0;
                15'h2FCC: d <= 8'hC0; 15'h2FCD: d <= 8'hC0; 15'h2FCE: d <= 8'hC0; 15'h2FCF: d <= 8'hC0;
                15'h2FD0: d <= 8'hC0; 15'h2FD1: d <= 8'hC0; 15'h2FD2: d <= 8'hC0; 15'h2FD3: d <= 8'hC0;
                15'h2FD4: d <= 8'hC0; 15'h2FD5: d <= 8'hC0; 15'h2FD6: d <= 8'hC0; 15'h2FD7: d <= 8'hC0;
                15'h2FD8: d <= 8'hC0; 15'h2FD9: d <= 8'hC0; 15'h2FDA: d <= 8'hC0; 15'h2FDB: d <= 8'hC0;
                15'h2FDC: d <= 8'hC0; 15'h2FDD: d <= 8'hC0; 15'h2FDE: d <= 8'hC0; 15'h2FDF: d <= 8'hC0;
                15'h2FE0: d <= 8'hC0; 15'h2FE1: d <= 8'hC0; 15'h2FE2: d <= 8'hC0; 15'h2FE3: d <= 8'hC0;
                15'h2FE4: d <= 8'hC0; 15'h2FE5: d <= 8'hC0; 15'h2FE6: d <= 8'hC0; 15'h2FE7: d <= 8'hC0;
                15'h2FE8: d <= 8'hC0; 15'h2FE9: d <= 8'hC0; 15'h2FEA: d <= 8'hC0; 15'h2FEB: d <= 8'hC0;
                15'h2FEC: d <= 8'hC0; 15'h2FED: d <= 8'hC0; 15'h2FEE: d <= 8'hC0; 15'h2FEF: d <= 8'hC0;
                15'h2FF0: d <= 8'hC0; 15'h2FF1: d <= 8'hC0; 15'h2FF2: d <= 8'hC0; 15'h2FF3: d <= 8'hC0;
                15'h2FF4: d <= 8'hC0; 15'h2FF5: d <= 8'hC0; 15'h2FF6: d <= 8'hC0; 15'h2FF7: d <= 8'hC0;
                15'h2FF8: d <= 8'hC0; 15'h2FF9: d <= 8'hC0; 15'h2FFA: d <= 8'hC0; 15'h2FFB: d <= 8'hC0;
                15'h2FFC: d <= 8'hC0; 15'h2FFD: d <= 8'hC0; 15'h2FFE: d <= 8'hC0; 15'h2FFF: d <= 8'hC0;
                15'h3000: d <= 8'hC0; 15'h3001: d <= 8'hC0; 15'h3002: d <= 8'hC0; 15'h3003: d <= 8'hC0;
                15'h3004: d <= 8'hC0; 15'h3005: d <= 8'hC0; 15'h3006: d <= 8'hC0; 15'h3007: d <= 8'hC0;
                15'h3008: d <= 8'hC0; 15'h3009: d <= 8'hC0; 15'h300A: d <= 8'hC0; 15'h300B: d <= 8'hC0;
                15'h300C: d <= 8'hC0; 15'h300D: d <= 8'hC0; 15'h300E: d <= 8'hC0; 15'h300F: d <= 8'hC0;
                15'h3010: d <= 8'hC0; 15'h3011: d <= 8'hC0; 15'h3012: d <= 8'hC0; 15'h3013: d <= 8'hC0;
                15'h3014: d <= 8'hC0; 15'h3015: d <= 8'hC0; 15'h3016: d <= 8'hC0; 15'h3017: d <= 8'hC0;
                15'h3018: d <= 8'hC0; 15'h3019: d <= 8'hC0; 15'h301A: d <= 8'hC0; 15'h301B: d <= 8'hC0;
                15'h301C: d <= 8'hC0; 15'h301D: d <= 8'hC0; 15'h301E: d <= 8'hC0; 15'h301F: d <= 8'hC0;
                15'h3020: d <= 8'hC0; 15'h3021: d <= 8'hC0; 15'h3022: d <= 8'hC0; 15'h3023: d <= 8'hC0;
                15'h3024: d <= 8'hC0; 15'h3025: d <= 8'hC0; 15'h3026: d <= 8'hC0; 15'h3027: d <= 8'hC0;
                15'h3028: d <= 8'hC0; 15'h3029: d <= 8'hC0; 15'h302A: d <= 8'hC0; 15'h302B: d <= 8'hC0;
                15'h302C: d <= 8'hC0; 15'h302D: d <= 8'hC0; 15'h302E: d <= 8'hC0; 15'h302F: d <= 8'hC0;
                15'h3030: d <= 8'hC0; 15'h3031: d <= 8'hC0; 15'h3032: d <= 8'hC0; 15'h3033: d <= 8'hC0;
                15'h3034: d <= 8'hC0; 15'h3035: d <= 8'hC0; 15'h3036: d <= 8'hC0; 15'h3037: d <= 8'hC0;
                15'h3038: d <= 8'hC0; 15'h3039: d <= 8'hC0; 15'h303A: d <= 8'hC0; 15'h303B: d <= 8'hC0;
                15'h303C: d <= 8'hC0; 15'h303D: d <= 8'hC0; 15'h303E: d <= 8'hC0; 15'h303F: d <= 8'hC0;
                15'h3040: d <= 8'hC0; 15'h3041: d <= 8'hC0; 15'h3042: d <= 8'hC0; 15'h3043: d <= 8'hC0;
                15'h3044: d <= 8'hC0; 15'h3045: d <= 8'hC0; 15'h3046: d <= 8'hC0; 15'h3047: d <= 8'hC0;
                15'h3048: d <= 8'hC0; 15'h3049: d <= 8'hC0; 15'h304A: d <= 8'hC0; 15'h304B: d <= 8'hC0;
                15'h304C: d <= 8'hC0; 15'h304D: d <= 8'hC0; 15'h304E: d <= 8'hC0; 15'h304F: d <= 8'hC0;
                15'h3050: d <= 8'hC0; 15'h3051: d <= 8'hC0; 15'h3052: d <= 8'hC0; 15'h3053: d <= 8'hC0;
                15'h3054: d <= 8'hC0; 15'h3055: d <= 8'hC0; 15'h3056: d <= 8'hC0; 15'h3057: d <= 8'hC0;
                15'h3058: d <= 8'hC0; 15'h3059: d <= 8'hC0; 15'h305A: d <= 8'hC0; 15'h305B: d <= 8'hC0;
                15'h305C: d <= 8'hC0; 15'h305D: d <= 8'hC0; 15'h305E: d <= 8'hC0; 15'h305F: d <= 8'hC0;
                15'h3060: d <= 8'hC0; 15'h3061: d <= 8'hC0; 15'h3062: d <= 8'hC0; 15'h3063: d <= 8'hC0;
                15'h3064: d <= 8'hC0; 15'h3065: d <= 8'hC0; 15'h3066: d <= 8'hC0; 15'h3067: d <= 8'hC0;
                15'h3068: d <= 8'hC0; 15'h3069: d <= 8'hC0; 15'h306A: d <= 8'hC0; 15'h306B: d <= 8'hC0;
                15'h306C: d <= 8'hC0; 15'h306D: d <= 8'hC0; 15'h306E: d <= 8'hC0; 15'h306F: d <= 8'hC0;
                15'h3070: d <= 8'hC0; 15'h3071: d <= 8'hC0; 15'h3072: d <= 8'hC0; 15'h3073: d <= 8'hC0;
                15'h3074: d <= 8'hC0; 15'h3075: d <= 8'hC0; 15'h3076: d <= 8'hC0; 15'h3077: d <= 8'hC0;
                15'h3078: d <= 8'hC0; 15'h3079: d <= 8'hC0; 15'h307A: d <= 8'hC0; 15'h307B: d <= 8'hC0;
                15'h307C: d <= 8'hC0; 15'h307D: d <= 8'hC0; 15'h307E: d <= 8'hC0; 15'h307F: d <= 8'hC0;
                15'h3080: d <= 8'hC0; 15'h3081: d <= 8'hC0; 15'h3082: d <= 8'hC0; 15'h3083: d <= 8'hC0;
                15'h3084: d <= 8'hC0; 15'h3085: d <= 8'hC0; 15'h3086: d <= 8'hC0; 15'h3087: d <= 8'hC0;
                15'h3088: d <= 8'hC0; 15'h3089: d <= 8'hC0; 15'h308A: d <= 8'hC0; 15'h308B: d <= 8'hC0;
                15'h308C: d <= 8'hC0; 15'h308D: d <= 8'hC0; 15'h308E: d <= 8'hC0; 15'h308F: d <= 8'hC0;
                15'h3090: d <= 8'hC0; 15'h3091: d <= 8'hC0; 15'h3092: d <= 8'hC0; 15'h3093: d <= 8'hC0;
                15'h3094: d <= 8'hC0; 15'h3095: d <= 8'hC0; 15'h3096: d <= 8'hC0; 15'h3097: d <= 8'hC0;
                15'h3098: d <= 8'hC0; 15'h3099: d <= 8'hC0; 15'h309A: d <= 8'hC0; 15'h309B: d <= 8'hC0;
                15'h309C: d <= 8'hC0; 15'h309D: d <= 8'hC0; 15'h309E: d <= 8'hC0; 15'h309F: d <= 8'hC0;
                15'h30A0: d <= 8'hC0; 15'h30A1: d <= 8'hC0; 15'h30A2: d <= 8'hC0; 15'h30A3: d <= 8'hC0;
                15'h30A4: d <= 8'hC0; 15'h30A5: d <= 8'hC0; 15'h30A6: d <= 8'hC0; 15'h30A7: d <= 8'hC0;
                15'h30A8: d <= 8'hC0; 15'h30A9: d <= 8'hC0; 15'h30AA: d <= 8'hC0; 15'h30AB: d <= 8'hC0;
                15'h30AC: d <= 8'hC0; 15'h30AD: d <= 8'hC0; 15'h30AE: d <= 8'hC0; 15'h30AF: d <= 8'hC0;
                15'h30B0: d <= 8'hC0; 15'h30B1: d <= 8'hC0; 15'h30B2: d <= 8'hC0; 15'h30B3: d <= 8'hC0;
                15'h30B4: d <= 8'hC0; 15'h30B5: d <= 8'hC0; 15'h30B6: d <= 8'hC0; 15'h30B7: d <= 8'hC0;
                15'h30B8: d <= 8'hC0; 15'h30B9: d <= 8'hC0; 15'h30BA: d <= 8'hC0; 15'h30BB: d <= 8'hC0;
                15'h30BC: d <= 8'hC0; 15'h30BD: d <= 8'hC0; 15'h30BE: d <= 8'hC0; 15'h30BF: d <= 8'hC0;
                15'h30C0: d <= 8'hC0; 15'h30C1: d <= 8'hC0; 15'h30C2: d <= 8'hC0; 15'h30C3: d <= 8'hC0;
                15'h30C4: d <= 8'hC0; 15'h30C5: d <= 8'hC0; 15'h30C6: d <= 8'hC0; 15'h30C7: d <= 8'hC0;
                15'h30C8: d <= 8'hC0; 15'h30C9: d <= 8'hC0; 15'h30CA: d <= 8'hC0; 15'h30CB: d <= 8'hC0;
                15'h30CC: d <= 8'hC0; 15'h30CD: d <= 8'hC0; 15'h30CE: d <= 8'hC0; 15'h30CF: d <= 8'hC0;
                15'h30D0: d <= 8'hC0; 15'h30D1: d <= 8'hC0; 15'h30D2: d <= 8'hC0; 15'h30D3: d <= 8'hC0;
                15'h30D4: d <= 8'hC0; 15'h30D5: d <= 8'hC0; 15'h30D6: d <= 8'hC0; 15'h30D7: d <= 8'hC0;
                15'h30D8: d <= 8'hC0; 15'h30D9: d <= 8'hC0; 15'h30DA: d <= 8'hC0; 15'h30DB: d <= 8'hC0;
                15'h30DC: d <= 8'hC0; 15'h30DD: d <= 8'hC0; 15'h30DE: d <= 8'hC0; 15'h30DF: d <= 8'hC0;
                15'h30E0: d <= 8'hC0; 15'h30E1: d <= 8'hC0; 15'h30E2: d <= 8'hC0; 15'h30E3: d <= 8'hC0;
                15'h30E4: d <= 8'hC0; 15'h30E5: d <= 8'hC0; 15'h30E6: d <= 8'hC0; 15'h30E7: d <= 8'hC0;
                15'h30E8: d <= 8'hC0; 15'h30E9: d <= 8'hC0; 15'h30EA: d <= 8'hC0; 15'h30EB: d <= 8'hC0;
                15'h30EC: d <= 8'hC0; 15'h30ED: d <= 8'hC0; 15'h30EE: d <= 8'hC0; 15'h30EF: d <= 8'hC0;
                15'h30F0: d <= 8'hC0; 15'h30F1: d <= 8'hC0; 15'h30F2: d <= 8'hC0; 15'h30F3: d <= 8'hC0;
                15'h30F4: d <= 8'hC0; 15'h30F5: d <= 8'hC0; 15'h30F6: d <= 8'hC0; 15'h30F7: d <= 8'hC0;
                15'h30F8: d <= 8'hC0; 15'h30F9: d <= 8'hC0; 15'h30FA: d <= 8'hC0; 15'h30FB: d <= 8'hC0;
                15'h30FC: d <= 8'hC0; 15'h30FD: d <= 8'hC0; 15'h30FE: d <= 8'hC0; 15'h30FF: d <= 8'hC0;
                15'h3100: d <= 8'hC0; 15'h3101: d <= 8'hC0; 15'h3102: d <= 8'hC0; 15'h3103: d <= 8'hC0;
                15'h3104: d <= 8'hC0; 15'h3105: d <= 8'hC0; 15'h3106: d <= 8'hC0; 15'h3107: d <= 8'hC0;
                15'h3108: d <= 8'hC0; 15'h3109: d <= 8'hC0; 15'h310A: d <= 8'hC0; 15'h310B: d <= 8'hC0;
                15'h310C: d <= 8'hC0; 15'h310D: d <= 8'hC0; 15'h310E: d <= 8'hC0; 15'h310F: d <= 8'hC0;
                15'h3110: d <= 8'hC0; 15'h3111: d <= 8'hC0; 15'h3112: d <= 8'hC0; 15'h3113: d <= 8'hC0;
                15'h3114: d <= 8'hC0; 15'h3115: d <= 8'hC0; 15'h3116: d <= 8'hC0; 15'h3117: d <= 8'hC0;
                15'h3118: d <= 8'hC0; 15'h3119: d <= 8'hC0; 15'h311A: d <= 8'hC0; 15'h311B: d <= 8'hC0;
                15'h311C: d <= 8'hC0; 15'h311D: d <= 8'hC0; 15'h311E: d <= 8'hC0; 15'h311F: d <= 8'hC0;
                15'h3120: d <= 8'hC0; 15'h3121: d <= 8'hC0; 15'h3122: d <= 8'hC0; 15'h3123: d <= 8'hC0;
                15'h3124: d <= 8'hC0; 15'h3125: d <= 8'hC0; 15'h3126: d <= 8'hC0; 15'h3127: d <= 8'hC0;
                15'h3128: d <= 8'hC0; 15'h3129: d <= 8'hC0; 15'h312A: d <= 8'hC0; 15'h312B: d <= 8'hC0;
                15'h312C: d <= 8'hC0; 15'h312D: d <= 8'hC0; 15'h312E: d <= 8'hC0; 15'h312F: d <= 8'hC0;
                15'h3130: d <= 8'hC0; 15'h3131: d <= 8'hC0; 15'h3132: d <= 8'hC0; 15'h3133: d <= 8'hC0;
                15'h3134: d <= 8'hC0; 15'h3135: d <= 8'hC0; 15'h3136: d <= 8'hC0; 15'h3137: d <= 8'hC0;
                15'h3138: d <= 8'hC0; 15'h3139: d <= 8'hC0; 15'h313A: d <= 8'hC0; 15'h313B: d <= 8'hC0;
                15'h313C: d <= 8'hC0; 15'h313D: d <= 8'hC0; 15'h313E: d <= 8'hC0; 15'h313F: d <= 8'hC0;
                15'h3140: d <= 8'hC0; 15'h3141: d <= 8'hC0; 15'h3142: d <= 8'hC0; 15'h3143: d <= 8'hC0;
                15'h3144: d <= 8'hC0; 15'h3145: d <= 8'hC0; 15'h3146: d <= 8'hC0; 15'h3147: d <= 8'hC0;
                15'h3148: d <= 8'hC0; 15'h3149: d <= 8'hC0; 15'h314A: d <= 8'hC0; 15'h314B: d <= 8'hC0;
                15'h314C: d <= 8'hC0; 15'h314D: d <= 8'hC0; 15'h314E: d <= 8'hC0; 15'h314F: d <= 8'hC0;
                15'h3150: d <= 8'hC0; 15'h3151: d <= 8'hC0; 15'h3152: d <= 8'hC0; 15'h3153: d <= 8'hC0;
                15'h3154: d <= 8'hC0; 15'h3155: d <= 8'hC0; 15'h3156: d <= 8'hC0; 15'h3157: d <= 8'hC0;
                15'h3158: d <= 8'hC0; 15'h3159: d <= 8'hC0; 15'h315A: d <= 8'hC0; 15'h315B: d <= 8'hC0;
                15'h315C: d <= 8'hC0; 15'h315D: d <= 8'hC0; 15'h315E: d <= 8'hC0; 15'h315F: d <= 8'hC0;
                15'h3160: d <= 8'hC0; 15'h3161: d <= 8'hC0; 15'h3162: d <= 8'hC0; 15'h3163: d <= 8'hC0;
                15'h3164: d <= 8'hC0; 15'h3165: d <= 8'hC0; 15'h3166: d <= 8'hC0; 15'h3167: d <= 8'hC0;
                15'h3168: d <= 8'hC0; 15'h3169: d <= 8'hC0; 15'h316A: d <= 8'hC0; 15'h316B: d <= 8'hC0;
                15'h316C: d <= 8'hC0; 15'h316D: d <= 8'hC0; 15'h316E: d <= 8'hC0; 15'h316F: d <= 8'hC0;
                15'h3170: d <= 8'hC0; 15'h3171: d <= 8'hC0; 15'h3172: d <= 8'hC0; 15'h3173: d <= 8'hC0;
                15'h3174: d <= 8'hC0; 15'h3175: d <= 8'hC0; 15'h3176: d <= 8'hC0; 15'h3177: d <= 8'hC0;
                15'h3178: d <= 8'hC0; 15'h3179: d <= 8'hC0; 15'h317A: d <= 8'hC0; 15'h317B: d <= 8'hC0;
                15'h317C: d <= 8'hC0; 15'h317D: d <= 8'hC0; 15'h317E: d <= 8'hC0; 15'h317F: d <= 8'hC0;
                15'h3180: d <= 8'hC0; 15'h3181: d <= 8'hC0; 15'h3182: d <= 8'hC0; 15'h3183: d <= 8'hC0;
                15'h3184: d <= 8'hC0; 15'h3185: d <= 8'hC0; 15'h3186: d <= 8'hC0; 15'h3187: d <= 8'hC0;
                15'h3188: d <= 8'hC0; 15'h3189: d <= 8'hC0; 15'h318A: d <= 8'hC0; 15'h318B: d <= 8'hC0;
                15'h318C: d <= 8'hC0; 15'h318D: d <= 8'hC0; 15'h318E: d <= 8'hC0; 15'h318F: d <= 8'hC0;
                15'h3190: d <= 8'hC0; 15'h3191: d <= 8'hC0; 15'h3192: d <= 8'hC0; 15'h3193: d <= 8'hC0;
                15'h3194: d <= 8'hC0; 15'h3195: d <= 8'hC0; 15'h3196: d <= 8'hC0; 15'h3197: d <= 8'hC0;
                15'h3198: d <= 8'hC0; 15'h3199: d <= 8'hC0; 15'h319A: d <= 8'hC0; 15'h319B: d <= 8'hC0;
                15'h319C: d <= 8'hC0; 15'h319D: d <= 8'hC0; 15'h319E: d <= 8'hC0; 15'h319F: d <= 8'hC0;
                15'h31A0: d <= 8'hC0; 15'h31A1: d <= 8'hC0; 15'h31A2: d <= 8'hC0; 15'h31A3: d <= 8'hC0;
                15'h31A4: d <= 8'hC0; 15'h31A5: d <= 8'hC0; 15'h31A6: d <= 8'hC0; 15'h31A7: d <= 8'hC0;
                15'h31A8: d <= 8'hC0; 15'h31A9: d <= 8'hC0; 15'h31AA: d <= 8'hC0; 15'h31AB: d <= 8'hC0;
                15'h31AC: d <= 8'hC0; 15'h31AD: d <= 8'hC0; 15'h31AE: d <= 8'hC0; 15'h31AF: d <= 8'hC0;
                15'h31B0: d <= 8'hC0; 15'h31B1: d <= 8'hC0; 15'h31B2: d <= 8'hC0; 15'h31B3: d <= 8'hC0;
                15'h31B4: d <= 8'hC0; 15'h31B5: d <= 8'hC0; 15'h31B6: d <= 8'hC0; 15'h31B7: d <= 8'hC0;
                15'h31B8: d <= 8'hC0; 15'h31B9: d <= 8'hC0; 15'h31BA: d <= 8'hC0; 15'h31BB: d <= 8'hC0;
                15'h31BC: d <= 8'hC0; 15'h31BD: d <= 8'hC0; 15'h31BE: d <= 8'hC0; 15'h31BF: d <= 8'hC0;
                15'h31C0: d <= 8'hC0; 15'h31C1: d <= 8'hC0; 15'h31C2: d <= 8'hC0; 15'h31C3: d <= 8'hC0;
                15'h31C4: d <= 8'hC0; 15'h31C5: d <= 8'hC0; 15'h31C6: d <= 8'hC0; 15'h31C7: d <= 8'hC0;
                15'h31C8: d <= 8'hC0; 15'h31C9: d <= 8'hC0; 15'h31CA: d <= 8'hC0; 15'h31CB: d <= 8'hC0;
                15'h31CC: d <= 8'hC0; 15'h31CD: d <= 8'hC0; 15'h31CE: d <= 8'hC0; 15'h31CF: d <= 8'hC0;
                15'h31D0: d <= 8'hC0; 15'h31D1: d <= 8'hC0; 15'h31D2: d <= 8'hC0; 15'h31D3: d <= 8'hC0;
                15'h31D4: d <= 8'hC0; 15'h31D5: d <= 8'hC0; 15'h31D6: d <= 8'hC0; 15'h31D7: d <= 8'hC0;
                15'h31D8: d <= 8'hC0; 15'h31D9: d <= 8'hC0; 15'h31DA: d <= 8'hC0; 15'h31DB: d <= 8'hC0;
                15'h31DC: d <= 8'hC0; 15'h31DD: d <= 8'hC0; 15'h31DE: d <= 8'hC0; 15'h31DF: d <= 8'hC0;
                15'h31E0: d <= 8'hC0; 15'h31E1: d <= 8'hC0; 15'h31E2: d <= 8'hC0; 15'h31E3: d <= 8'hC0;
                15'h31E4: d <= 8'hC0; 15'h31E5: d <= 8'hC0; 15'h31E6: d <= 8'hC0; 15'h31E7: d <= 8'hC0;
                15'h31E8: d <= 8'hC0; 15'h31E9: d <= 8'hC0; 15'h31EA: d <= 8'hC0; 15'h31EB: d <= 8'hC0;
                15'h31EC: d <= 8'hC0; 15'h31ED: d <= 8'hC0; 15'h31EE: d <= 8'hC0; 15'h31EF: d <= 8'hC0;
                15'h31F0: d <= 8'hC0; 15'h31F1: d <= 8'hC0; 15'h31F2: d <= 8'hC0; 15'h31F3: d <= 8'hC0;
                15'h31F4: d <= 8'hC0; 15'h31F5: d <= 8'hC0; 15'h31F6: d <= 8'hC0; 15'h31F7: d <= 8'hC0;
                15'h31F8: d <= 8'hC0; 15'h31F9: d <= 8'hC0; 15'h31FA: d <= 8'hC0; 15'h31FB: d <= 8'hC0;
                15'h31FC: d <= 8'hC0; 15'h31FD: d <= 8'hC0; 15'h31FE: d <= 8'hC0; 15'h31FF: d <= 8'hC0;
                15'h3200: d <= 8'hC0; 15'h3201: d <= 8'hC0; 15'h3202: d <= 8'hC0; 15'h3203: d <= 8'hC0;
                15'h3204: d <= 8'hC0; 15'h3205: d <= 8'hC0; 15'h3206: d <= 8'hC0; 15'h3207: d <= 8'hC0;
                15'h3208: d <= 8'hC0; 15'h3209: d <= 8'hC0; 15'h320A: d <= 8'hC0; 15'h320B: d <= 8'hC0;
                15'h320C: d <= 8'hC0; 15'h320D: d <= 8'hC0; 15'h320E: d <= 8'hC0; 15'h320F: d <= 8'hC0;
                15'h3210: d <= 8'hC0; 15'h3211: d <= 8'hC0; 15'h3212: d <= 8'hC0; 15'h3213: d <= 8'hC0;
                15'h3214: d <= 8'hC0; 15'h3215: d <= 8'hC0; 15'h3216: d <= 8'hC0; 15'h3217: d <= 8'hC0;
                15'h3218: d <= 8'hC0; 15'h3219: d <= 8'hC0; 15'h321A: d <= 8'hC0; 15'h321B: d <= 8'hC0;
                15'h321C: d <= 8'hC0; 15'h321D: d <= 8'hC0; 15'h321E: d <= 8'hC0; 15'h321F: d <= 8'hC0;
                15'h3220: d <= 8'hC0; 15'h3221: d <= 8'hC0; 15'h3222: d <= 8'hC0; 15'h3223: d <= 8'hC0;
                15'h3224: d <= 8'hC0; 15'h3225: d <= 8'hC0; 15'h3226: d <= 8'hC0; 15'h3227: d <= 8'hC0;
                15'h3228: d <= 8'hC0; 15'h3229: d <= 8'hC0; 15'h322A: d <= 8'hC0; 15'h322B: d <= 8'hC0;
                15'h322C: d <= 8'hC0; 15'h322D: d <= 8'hC0; 15'h322E: d <= 8'hC0; 15'h322F: d <= 8'hC0;
                15'h3230: d <= 8'hC0; 15'h3231: d <= 8'hC0; 15'h3232: d <= 8'hC0; 15'h3233: d <= 8'hC0;
                15'h3234: d <= 8'hC0; 15'h3235: d <= 8'hC0; 15'h3236: d <= 8'hC0; 15'h3237: d <= 8'hC0;
                15'h3238: d <= 8'hC0; 15'h3239: d <= 8'hC0; 15'h323A: d <= 8'hC0; 15'h323B: d <= 8'hC0;
                15'h323C: d <= 8'hC0; 15'h323D: d <= 8'hC0; 15'h323E: d <= 8'hC0; 15'h323F: d <= 8'hC0;
                15'h3240: d <= 8'hC0; 15'h3241: d <= 8'hC0; 15'h3242: d <= 8'hC0; 15'h3243: d <= 8'hC0;
                15'h3244: d <= 8'hC0; 15'h3245: d <= 8'hC0; 15'h3246: d <= 8'hC0; 15'h3247: d <= 8'hC0;
                15'h3248: d <= 8'hC0; 15'h3249: d <= 8'hC0; 15'h324A: d <= 8'hC0; 15'h324B: d <= 8'hC0;
                15'h324C: d <= 8'hC0; 15'h324D: d <= 8'hC0; 15'h324E: d <= 8'hC0; 15'h324F: d <= 8'hC0;
                15'h3250: d <= 8'hC0; 15'h3251: d <= 8'hC0; 15'h3252: d <= 8'hC0; 15'h3253: d <= 8'hC0;
                15'h3254: d <= 8'hC0; 15'h3255: d <= 8'hC0; 15'h3256: d <= 8'hC0; 15'h3257: d <= 8'hC0;
                15'h3258: d <= 8'hC0; 15'h3259: d <= 8'hC0; 15'h325A: d <= 8'hC0; 15'h325B: d <= 8'hC0;
                15'h325C: d <= 8'hC0; 15'h325D: d <= 8'hC0; 15'h325E: d <= 8'hC0; 15'h325F: d <= 8'hC0;
                15'h3260: d <= 8'hC0; 15'h3261: d <= 8'hC0; 15'h3262: d <= 8'hC0; 15'h3263: d <= 8'hC0;
                15'h3264: d <= 8'hC0; 15'h3265: d <= 8'hC0; 15'h3266: d <= 8'hC0; 15'h3267: d <= 8'hC0;
                15'h3268: d <= 8'hC0; 15'h3269: d <= 8'hC0; 15'h326A: d <= 8'hC0; 15'h326B: d <= 8'hC0;
                15'h326C: d <= 8'hC0; 15'h326D: d <= 8'hC0; 15'h326E: d <= 8'hC0; 15'h326F: d <= 8'hC0;
                15'h3270: d <= 8'hC0; 15'h3271: d <= 8'hC0; 15'h3272: d <= 8'hC0; 15'h3273: d <= 8'hC0;
                15'h3274: d <= 8'hC0; 15'h3275: d <= 8'hC0; 15'h3276: d <= 8'hC0; 15'h3277: d <= 8'hC0;
                15'h3278: d <= 8'hC0; 15'h3279: d <= 8'hC0; 15'h327A: d <= 8'hC0; 15'h327B: d <= 8'hC0;
                15'h327C: d <= 8'hC0; 15'h327D: d <= 8'hC0; 15'h327E: d <= 8'hC0; 15'h327F: d <= 8'hC0;
                15'h3280: d <= 8'hC0; 15'h3281: d <= 8'hC0; 15'h3282: d <= 8'hC0; 15'h3283: d <= 8'hC0;
                15'h3284: d <= 8'hC0; 15'h3285: d <= 8'hC0; 15'h3286: d <= 8'hC0; 15'h3287: d <= 8'hC0;
                15'h3288: d <= 8'hC0; 15'h3289: d <= 8'hC0; 15'h328A: d <= 8'hC0; 15'h328B: d <= 8'hC0;
                15'h328C: d <= 8'hC0; 15'h328D: d <= 8'hC0; 15'h328E: d <= 8'hC0; 15'h328F: d <= 8'hC0;
                15'h3290: d <= 8'hC0; 15'h3291: d <= 8'hC0; 15'h3292: d <= 8'hC0; 15'h3293: d <= 8'hC0;
                15'h3294: d <= 8'hC0; 15'h3295: d <= 8'hC0; 15'h3296: d <= 8'hC0; 15'h3297: d <= 8'hC0;
                15'h3298: d <= 8'hC0; 15'h3299: d <= 8'hC0; 15'h329A: d <= 8'hC0; 15'h329B: d <= 8'hC0;
                15'h329C: d <= 8'hC0; 15'h329D: d <= 8'hC0; 15'h329E: d <= 8'hC0; 15'h329F: d <= 8'hC0;
                15'h32A0: d <= 8'hC0; 15'h32A1: d <= 8'hC0; 15'h32A2: d <= 8'hC0; 15'h32A3: d <= 8'hC0;
                15'h32A4: d <= 8'hC0; 15'h32A5: d <= 8'hC0; 15'h32A6: d <= 8'hC0; 15'h32A7: d <= 8'hC0;
                15'h32A8: d <= 8'hC0; 15'h32A9: d <= 8'hC0; 15'h32AA: d <= 8'hC0; 15'h32AB: d <= 8'hC0;
                15'h32AC: d <= 8'hC0; 15'h32AD: d <= 8'hC0; 15'h32AE: d <= 8'hC0; 15'h32AF: d <= 8'hC0;
                15'h32B0: d <= 8'hC0; 15'h32B1: d <= 8'hC0; 15'h32B2: d <= 8'hC0; 15'h32B3: d <= 8'hC0;
                15'h32B4: d <= 8'hC0; 15'h32B5: d <= 8'hC0; 15'h32B6: d <= 8'hC0; 15'h32B7: d <= 8'hC0;
                15'h32B8: d <= 8'hC0; 15'h32B9: d <= 8'hC0; 15'h32BA: d <= 8'hC0; 15'h32BB: d <= 8'hC0;
                15'h32BC: d <= 8'hC0; 15'h32BD: d <= 8'hC0; 15'h32BE: d <= 8'hC0; 15'h32BF: d <= 8'hC0;
                15'h32C0: d <= 8'hC0; 15'h32C1: d <= 8'hC0; 15'h32C2: d <= 8'hC0; 15'h32C3: d <= 8'hC0;
                15'h32C4: d <= 8'hC0; 15'h32C5: d <= 8'hC0; 15'h32C6: d <= 8'hC0; 15'h32C7: d <= 8'hC0;
                15'h32C8: d <= 8'hC0; 15'h32C9: d <= 8'hC0; 15'h32CA: d <= 8'hC0; 15'h32CB: d <= 8'hC0;
                15'h32CC: d <= 8'hC0; 15'h32CD: d <= 8'hC0; 15'h32CE: d <= 8'hC0; 15'h32CF: d <= 8'hC0;
                15'h32D0: d <= 8'hC0; 15'h32D1: d <= 8'hC0; 15'h32D2: d <= 8'hC0; 15'h32D3: d <= 8'hC0;
                15'h32D4: d <= 8'hC0; 15'h32D5: d <= 8'hC0; 15'h32D6: d <= 8'hC0; 15'h32D7: d <= 8'hC0;
                15'h32D8: d <= 8'hC0; 15'h32D9: d <= 8'hC0; 15'h32DA: d <= 8'hC0; 15'h32DB: d <= 8'hC0;
                15'h32DC: d <= 8'hC0; 15'h32DD: d <= 8'hC0; 15'h32DE: d <= 8'hC0; 15'h32DF: d <= 8'hC0;
                15'h32E0: d <= 8'hC0; 15'h32E1: d <= 8'hC0; 15'h32E2: d <= 8'hC0; 15'h32E3: d <= 8'hC0;
                15'h32E4: d <= 8'hC0; 15'h32E5: d <= 8'hC0; 15'h32E6: d <= 8'hC0; 15'h32E7: d <= 8'hC0;
                15'h32E8: d <= 8'hC0; 15'h32E9: d <= 8'hC0; 15'h32EA: d <= 8'hC0; 15'h32EB: d <= 8'hC0;
                15'h32EC: d <= 8'hC0; 15'h32ED: d <= 8'hC0; 15'h32EE: d <= 8'hC0; 15'h32EF: d <= 8'hC0;
                15'h32F0: d <= 8'hC0; 15'h32F1: d <= 8'hC0; 15'h32F2: d <= 8'hC0; 15'h32F3: d <= 8'hC0;
                15'h32F4: d <= 8'hC0; 15'h32F5: d <= 8'hC0; 15'h32F6: d <= 8'hC0; 15'h32F7: d <= 8'hC0;
                15'h32F8: d <= 8'hC0; 15'h32F9: d <= 8'hC0; 15'h32FA: d <= 8'hC0; 15'h32FB: d <= 8'hC0;
                15'h32FC: d <= 8'hC0; 15'h32FD: d <= 8'hC0; 15'h32FE: d <= 8'hC0; 15'h32FF: d <= 8'hC0;
                15'h3300: d <= 8'hC0; 15'h3301: d <= 8'hC0; 15'h3302: d <= 8'hC0; 15'h3303: d <= 8'hC0;
                15'h3304: d <= 8'hC0; 15'h3305: d <= 8'hC0; 15'h3306: d <= 8'hC0; 15'h3307: d <= 8'hC0;
                15'h3308: d <= 8'hC0; 15'h3309: d <= 8'hC0; 15'h330A: d <= 8'hC0; 15'h330B: d <= 8'hC0;
                15'h330C: d <= 8'hC0; 15'h330D: d <= 8'hC0; 15'h330E: d <= 8'hC0; 15'h330F: d <= 8'hC0;
                15'h3310: d <= 8'hC0; 15'h3311: d <= 8'hC0; 15'h3312: d <= 8'hC0; 15'h3313: d <= 8'hC0;
                15'h3314: d <= 8'hC0; 15'h3315: d <= 8'hC0; 15'h3316: d <= 8'hC0; 15'h3317: d <= 8'hC0;
                15'h3318: d <= 8'hC0; 15'h3319: d <= 8'hC0; 15'h331A: d <= 8'hC0; 15'h331B: d <= 8'hC0;
                15'h331C: d <= 8'hC0; 15'h331D: d <= 8'hC0; 15'h331E: d <= 8'hC0; 15'h331F: d <= 8'hC0;
                15'h3320: d <= 8'hC0; 15'h3321: d <= 8'hC0; 15'h3322: d <= 8'hC0; 15'h3323: d <= 8'hC0;
                15'h3324: d <= 8'hC0; 15'h3325: d <= 8'hC0; 15'h3326: d <= 8'hC0; 15'h3327: d <= 8'hC0;
                15'h3328: d <= 8'hC0; 15'h3329: d <= 8'hC0; 15'h332A: d <= 8'hC0; 15'h332B: d <= 8'hC0;
                15'h332C: d <= 8'hC0; 15'h332D: d <= 8'hC0; 15'h332E: d <= 8'hC0; 15'h332F: d <= 8'hC0;
                15'h3330: d <= 8'hC0; 15'h3331: d <= 8'hC0; 15'h3332: d <= 8'hC0; 15'h3333: d <= 8'hC0;
                15'h3334: d <= 8'hC0; 15'h3335: d <= 8'hC0; 15'h3336: d <= 8'hC0; 15'h3337: d <= 8'hC0;
                15'h3338: d <= 8'hC0; 15'h3339: d <= 8'hC0; 15'h333A: d <= 8'hC0; 15'h333B: d <= 8'hC0;
                15'h333C: d <= 8'hC0; 15'h333D: d <= 8'hC0; 15'h333E: d <= 8'hC0; 15'h333F: d <= 8'hC0;
                15'h3340: d <= 8'hC0; 15'h3341: d <= 8'hC0; 15'h3342: d <= 8'hC0; 15'h3343: d <= 8'hC0;
                15'h3344: d <= 8'hC0; 15'h3345: d <= 8'hC0; 15'h3346: d <= 8'hC0; 15'h3347: d <= 8'hC0;
                15'h3348: d <= 8'hC0; 15'h3349: d <= 8'hC0; 15'h334A: d <= 8'hC0; 15'h334B: d <= 8'hC0;
                15'h334C: d <= 8'hC0; 15'h334D: d <= 8'hC0; 15'h334E: d <= 8'hC0; 15'h334F: d <= 8'hC0;
                15'h3350: d <= 8'hC0; 15'h3351: d <= 8'hC0; 15'h3352: d <= 8'hC0; 15'h3353: d <= 8'hC0;
                15'h3354: d <= 8'hC0; 15'h3355: d <= 8'hC0; 15'h3356: d <= 8'hC0; 15'h3357: d <= 8'hC0;
                15'h3358: d <= 8'hC0; 15'h3359: d <= 8'hC0; 15'h335A: d <= 8'hC0; 15'h335B: d <= 8'hC0;
                15'h335C: d <= 8'hC0; 15'h335D: d <= 8'hC0; 15'h335E: d <= 8'hC0; 15'h335F: d <= 8'hC0;
                15'h3360: d <= 8'hC0; 15'h3361: d <= 8'hC0; 15'h3362: d <= 8'hC0; 15'h3363: d <= 8'hC0;
                15'h3364: d <= 8'hC0; 15'h3365: d <= 8'hC0; 15'h3366: d <= 8'hC0; 15'h3367: d <= 8'hC0;
                15'h3368: d <= 8'hC0; 15'h3369: d <= 8'hC0; 15'h336A: d <= 8'hC0; 15'h336B: d <= 8'hC0;
                15'h336C: d <= 8'hC0; 15'h336D: d <= 8'hC0; 15'h336E: d <= 8'hC0; 15'h336F: d <= 8'hC0;
                15'h3370: d <= 8'hC0; 15'h3371: d <= 8'hC0; 15'h3372: d <= 8'hC0; 15'h3373: d <= 8'hC0;
                15'h3374: d <= 8'hC0; 15'h3375: d <= 8'hC0; 15'h3376: d <= 8'hC0; 15'h3377: d <= 8'hC0;
                15'h3378: d <= 8'hC0; 15'h3379: d <= 8'hC0; 15'h337A: d <= 8'hC0; 15'h337B: d <= 8'hC0;
                15'h337C: d <= 8'hC0; 15'h337D: d <= 8'hC0; 15'h337E: d <= 8'hC0; 15'h337F: d <= 8'hC0;
                15'h3380: d <= 8'hC0; 15'h3381: d <= 8'hC0; 15'h3382: d <= 8'hC0; 15'h3383: d <= 8'hC0;
                15'h3384: d <= 8'hC0; 15'h3385: d <= 8'hC0; 15'h3386: d <= 8'hC0; 15'h3387: d <= 8'hC0;
                15'h3388: d <= 8'hC0; 15'h3389: d <= 8'hC0; 15'h338A: d <= 8'hC0; 15'h338B: d <= 8'hC0;
                15'h338C: d <= 8'hC0; 15'h338D: d <= 8'hC0; 15'h338E: d <= 8'hC0; 15'h338F: d <= 8'hC0;
                15'h3390: d <= 8'hC0; 15'h3391: d <= 8'hC0; 15'h3392: d <= 8'hC0; 15'h3393: d <= 8'hC0;
                15'h3394: d <= 8'hC0; 15'h3395: d <= 8'hC0; 15'h3396: d <= 8'hC0; 15'h3397: d <= 8'hC0;
                15'h3398: d <= 8'hC0; 15'h3399: d <= 8'hC0; 15'h339A: d <= 8'hC0; 15'h339B: d <= 8'hC0;
                15'h339C: d <= 8'hC0; 15'h339D: d <= 8'hC0; 15'h339E: d <= 8'hC0; 15'h339F: d <= 8'hC0;
                15'h33A0: d <= 8'hC0; 15'h33A1: d <= 8'hC0; 15'h33A2: d <= 8'hC0; 15'h33A3: d <= 8'hC0;
                15'h33A4: d <= 8'hC0; 15'h33A5: d <= 8'hC0; 15'h33A6: d <= 8'hC0; 15'h33A7: d <= 8'hC0;
                15'h33A8: d <= 8'hC0; 15'h33A9: d <= 8'hC0; 15'h33AA: d <= 8'hC0; 15'h33AB: d <= 8'hC0;
                15'h33AC: d <= 8'hC0; 15'h33AD: d <= 8'hC0; 15'h33AE: d <= 8'hC0; 15'h33AF: d <= 8'hC0;
                15'h33B0: d <= 8'hC0; 15'h33B1: d <= 8'hC0; 15'h33B2: d <= 8'hC0; 15'h33B3: d <= 8'hC0;
                15'h33B4: d <= 8'hC0; 15'h33B5: d <= 8'hC0; 15'h33B6: d <= 8'hC0; 15'h33B7: d <= 8'hC0;
                15'h33B8: d <= 8'hC0; 15'h33B9: d <= 8'hC0; 15'h33BA: d <= 8'hC0; 15'h33BB: d <= 8'hC0;
                15'h33BC: d <= 8'hC0; 15'h33BD: d <= 8'hC0; 15'h33BE: d <= 8'hC0; 15'h33BF: d <= 8'hC0;
                15'h33C0: d <= 8'hC0; 15'h33C1: d <= 8'hC0; 15'h33C2: d <= 8'hC0; 15'h33C3: d <= 8'hC0;
                15'h33C4: d <= 8'hC0; 15'h33C5: d <= 8'hC0; 15'h33C6: d <= 8'hC0; 15'h33C7: d <= 8'hC0;
                15'h33C8: d <= 8'hC0; 15'h33C9: d <= 8'hC0; 15'h33CA: d <= 8'hC0; 15'h33CB: d <= 8'hC0;
                15'h33CC: d <= 8'hC0; 15'h33CD: d <= 8'hC0; 15'h33CE: d <= 8'hC0; 15'h33CF: d <= 8'hC0;
                15'h33D0: d <= 8'hC0; 15'h33D1: d <= 8'hC0; 15'h33D2: d <= 8'hC0; 15'h33D3: d <= 8'hC0;
                15'h33D4: d <= 8'hC0; 15'h33D5: d <= 8'hC0; 15'h33D6: d <= 8'hC0; 15'h33D7: d <= 8'hC0;
                15'h33D8: d <= 8'hC0; 15'h33D9: d <= 8'hC0; 15'h33DA: d <= 8'hC0; 15'h33DB: d <= 8'hC0;
                15'h33DC: d <= 8'hC0; 15'h33DD: d <= 8'hC0; 15'h33DE: d <= 8'hC0; 15'h33DF: d <= 8'hC0;
                15'h33E0: d <= 8'hC0; 15'h33E1: d <= 8'hC0; 15'h33E2: d <= 8'hC0; 15'h33E3: d <= 8'hC0;
                15'h33E4: d <= 8'hC0; 15'h33E5: d <= 8'hC0; 15'h33E6: d <= 8'hC0; 15'h33E7: d <= 8'hC0;
                15'h33E8: d <= 8'hC0; 15'h33E9: d <= 8'hC0; 15'h33EA: d <= 8'hC0; 15'h33EB: d <= 8'hC0;
                15'h33EC: d <= 8'hC0; 15'h33ED: d <= 8'hC0; 15'h33EE: d <= 8'hC0; 15'h33EF: d <= 8'hC0;
                15'h33F0: d <= 8'hC0; 15'h33F1: d <= 8'hC0; 15'h33F2: d <= 8'hC0; 15'h33F3: d <= 8'hC0;
                15'h33F4: d <= 8'hC0; 15'h33F5: d <= 8'hC0; 15'h33F6: d <= 8'hC0; 15'h33F7: d <= 8'hC0;
                15'h33F8: d <= 8'hC0; 15'h33F9: d <= 8'hC0; 15'h33FA: d <= 8'hC0; 15'h33FB: d <= 8'hC0;
                15'h33FC: d <= 8'hC0; 15'h33FD: d <= 8'hC0; 15'h33FE: d <= 8'hC0; 15'h33FF: d <= 8'hC0;
                15'h3400: d <= 8'hC0; 15'h3401: d <= 8'hC0; 15'h3402: d <= 8'hC0; 15'h3403: d <= 8'hC0;
                15'h3404: d <= 8'hC0; 15'h3405: d <= 8'hC0; 15'h3406: d <= 8'hC0; 15'h3407: d <= 8'hC0;
                15'h3408: d <= 8'hC0; 15'h3409: d <= 8'hC0; 15'h340A: d <= 8'hC0; 15'h340B: d <= 8'hC0;
                15'h340C: d <= 8'hC0; 15'h340D: d <= 8'hC0; 15'h340E: d <= 8'hC0; 15'h340F: d <= 8'hC0;
                15'h3410: d <= 8'hC0; 15'h3411: d <= 8'hC0; 15'h3412: d <= 8'hC0; 15'h3413: d <= 8'hC0;
                15'h3414: d <= 8'hC0; 15'h3415: d <= 8'hC0; 15'h3416: d <= 8'hC0; 15'h3417: d <= 8'hC0;
                15'h3418: d <= 8'hC0; 15'h3419: d <= 8'hC0; 15'h341A: d <= 8'hC0; 15'h341B: d <= 8'hC0;
                15'h341C: d <= 8'hC0; 15'h341D: d <= 8'hC0; 15'h341E: d <= 8'hC0; 15'h341F: d <= 8'hC0;
                15'h3420: d <= 8'hC0; 15'h3421: d <= 8'hC0; 15'h3422: d <= 8'hC0; 15'h3423: d <= 8'hC0;
                15'h3424: d <= 8'hC0; 15'h3425: d <= 8'hC0; 15'h3426: d <= 8'hC0; 15'h3427: d <= 8'hC0;
                15'h3428: d <= 8'hC0; 15'h3429: d <= 8'hC0; 15'h342A: d <= 8'hC0; 15'h342B: d <= 8'hC0;
                15'h342C: d <= 8'hC0; 15'h342D: d <= 8'hC0; 15'h342E: d <= 8'hC0; 15'h342F: d <= 8'hC0;
                15'h3430: d <= 8'hC0; 15'h3431: d <= 8'hC0; 15'h3432: d <= 8'hC0; 15'h3433: d <= 8'hC0;
                15'h3434: d <= 8'hC0; 15'h3435: d <= 8'hC0; 15'h3436: d <= 8'hC0; 15'h3437: d <= 8'hC0;
                15'h3438: d <= 8'hC0; 15'h3439: d <= 8'hC0; 15'h343A: d <= 8'hC0; 15'h343B: d <= 8'hC0;
                15'h343C: d <= 8'hC0; 15'h343D: d <= 8'hC0; 15'h343E: d <= 8'hC0; 15'h343F: d <= 8'hC0;
                15'h3440: d <= 8'hC0; 15'h3441: d <= 8'hC0; 15'h3442: d <= 8'hC0; 15'h3443: d <= 8'hC0;
                15'h3444: d <= 8'hC0; 15'h3445: d <= 8'hC0; 15'h3446: d <= 8'hC0; 15'h3447: d <= 8'hC0;
                15'h3448: d <= 8'hC0; 15'h3449: d <= 8'hC0; 15'h344A: d <= 8'hC0; 15'h344B: d <= 8'hC0;
                15'h344C: d <= 8'hC0; 15'h344D: d <= 8'hC0; 15'h344E: d <= 8'hC0; 15'h344F: d <= 8'hC0;
                15'h3450: d <= 8'hC0; 15'h3451: d <= 8'hC0; 15'h3452: d <= 8'hC0; 15'h3453: d <= 8'hC0;
                15'h3454: d <= 8'hC0; 15'h3455: d <= 8'hC0; 15'h3456: d <= 8'hC0; 15'h3457: d <= 8'hC0;
                15'h3458: d <= 8'hC0; 15'h3459: d <= 8'hC0; 15'h345A: d <= 8'hC0; 15'h345B: d <= 8'hC0;
                15'h345C: d <= 8'hC0; 15'h345D: d <= 8'hC0; 15'h345E: d <= 8'hC0; 15'h345F: d <= 8'hC0;
                15'h3460: d <= 8'hC0; 15'h3461: d <= 8'hC0; 15'h3462: d <= 8'hC0; 15'h3463: d <= 8'hC0;
                15'h3464: d <= 8'hC0; 15'h3465: d <= 8'hC0; 15'h3466: d <= 8'hC0; 15'h3467: d <= 8'hC0;
                15'h3468: d <= 8'hC0; 15'h3469: d <= 8'hC0; 15'h346A: d <= 8'hC0; 15'h346B: d <= 8'hC0;
                15'h346C: d <= 8'hC0; 15'h346D: d <= 8'hC0; 15'h346E: d <= 8'hC0; 15'h346F: d <= 8'hC0;
                15'h3470: d <= 8'hC0; 15'h3471: d <= 8'hC0; 15'h3472: d <= 8'hC0; 15'h3473: d <= 8'hC0;
                15'h3474: d <= 8'hC0; 15'h3475: d <= 8'hC0; 15'h3476: d <= 8'hC0; 15'h3477: d <= 8'hC0;
                15'h3478: d <= 8'hC0; 15'h3479: d <= 8'hC0; 15'h347A: d <= 8'hC0; 15'h347B: d <= 8'hC0;
                15'h347C: d <= 8'hC0; 15'h347D: d <= 8'hC0; 15'h347E: d <= 8'hC0; 15'h347F: d <= 8'hC0;
                15'h3480: d <= 8'hC0; 15'h3481: d <= 8'hC0; 15'h3482: d <= 8'hC0; 15'h3483: d <= 8'hC0;
                15'h3484: d <= 8'hC0; 15'h3485: d <= 8'hC0; 15'h3486: d <= 8'hC0; 15'h3487: d <= 8'hC0;
                15'h3488: d <= 8'hC0; 15'h3489: d <= 8'hC0; 15'h348A: d <= 8'hC0; 15'h348B: d <= 8'hC0;
                15'h348C: d <= 8'hC0; 15'h348D: d <= 8'hC0; 15'h348E: d <= 8'hC0; 15'h348F: d <= 8'hC0;
                15'h3490: d <= 8'hC0; 15'h3491: d <= 8'hC0; 15'h3492: d <= 8'hC0; 15'h3493: d <= 8'hC0;
                15'h3494: d <= 8'hC0; 15'h3495: d <= 8'hC0; 15'h3496: d <= 8'hC0; 15'h3497: d <= 8'hC0;
                15'h3498: d <= 8'hC0; 15'h3499: d <= 8'hC0; 15'h349A: d <= 8'hC0; 15'h349B: d <= 8'hC0;
                15'h349C: d <= 8'hC0; 15'h349D: d <= 8'hC0; 15'h349E: d <= 8'hC0; 15'h349F: d <= 8'hC0;
                15'h34A0: d <= 8'hC0; 15'h34A1: d <= 8'hC0; 15'h34A2: d <= 8'hC0; 15'h34A3: d <= 8'hC0;
                15'h34A4: d <= 8'hC0; 15'h34A5: d <= 8'hC0; 15'h34A6: d <= 8'hC0; 15'h34A7: d <= 8'hC0;
                15'h34A8: d <= 8'hC0; 15'h34A9: d <= 8'hC0; 15'h34AA: d <= 8'hC0; 15'h34AB: d <= 8'hC0;
                15'h34AC: d <= 8'hC0; 15'h34AD: d <= 8'hC0; 15'h34AE: d <= 8'hC0; 15'h34AF: d <= 8'hC0;
                15'h34B0: d <= 8'hC0; 15'h34B1: d <= 8'hC0; 15'h34B2: d <= 8'hC0; 15'h34B3: d <= 8'hC0;
                15'h34B4: d <= 8'hC0; 15'h34B5: d <= 8'hC0; 15'h34B6: d <= 8'hC0; 15'h34B7: d <= 8'hC0;
                15'h34B8: d <= 8'hC0; 15'h34B9: d <= 8'hC0; 15'h34BA: d <= 8'hC0; 15'h34BB: d <= 8'hC0;
                15'h34BC: d <= 8'hC0; 15'h34BD: d <= 8'hC0; 15'h34BE: d <= 8'hC0; 15'h34BF: d <= 8'hC0;
                15'h34C0: d <= 8'hC0; 15'h34C1: d <= 8'hC0; 15'h34C2: d <= 8'hC0; 15'h34C3: d <= 8'hC0;
                15'h34C4: d <= 8'hC0; 15'h34C5: d <= 8'hC0; 15'h34C6: d <= 8'hC0; 15'h34C7: d <= 8'hC0;
                15'h34C8: d <= 8'hC0; 15'h34C9: d <= 8'hC0; 15'h34CA: d <= 8'hC0; 15'h34CB: d <= 8'hC0;
                15'h34CC: d <= 8'hC0; 15'h34CD: d <= 8'hC0; 15'h34CE: d <= 8'hC0; 15'h34CF: d <= 8'hC0;
                15'h34D0: d <= 8'hC0; 15'h34D1: d <= 8'hC0; 15'h34D2: d <= 8'hC0; 15'h34D3: d <= 8'hC0;
                15'h34D4: d <= 8'hC0; 15'h34D5: d <= 8'hC0; 15'h34D6: d <= 8'hC0; 15'h34D7: d <= 8'hC0;
                15'h34D8: d <= 8'hC0; 15'h34D9: d <= 8'hC0; 15'h34DA: d <= 8'hC0; 15'h34DB: d <= 8'hC0;
                15'h34DC: d <= 8'hC0; 15'h34DD: d <= 8'hC0; 15'h34DE: d <= 8'hC0; 15'h34DF: d <= 8'hC0;
                15'h34E0: d <= 8'hC0; 15'h34E1: d <= 8'hC0; 15'h34E2: d <= 8'hC0; 15'h34E3: d <= 8'hC0;
                15'h34E4: d <= 8'hC0; 15'h34E5: d <= 8'hC0; 15'h34E6: d <= 8'hC0; 15'h34E7: d <= 8'hC0;
                15'h34E8: d <= 8'hC0; 15'h34E9: d <= 8'hC0; 15'h34EA: d <= 8'hC0; 15'h34EB: d <= 8'hC0;
                15'h34EC: d <= 8'hC0; 15'h34ED: d <= 8'hC0; 15'h34EE: d <= 8'hC0; 15'h34EF: d <= 8'hC0;
                15'h34F0: d <= 8'hC0; 15'h34F1: d <= 8'hC0; 15'h34F2: d <= 8'hC0; 15'h34F3: d <= 8'hC0;
                15'h34F4: d <= 8'hC0; 15'h34F5: d <= 8'hC0; 15'h34F6: d <= 8'hC0; 15'h34F7: d <= 8'hC0;
                15'h34F8: d <= 8'hC0; 15'h34F9: d <= 8'hC0; 15'h34FA: d <= 8'hC0; 15'h34FB: d <= 8'hC0;
                15'h34FC: d <= 8'hC0; 15'h34FD: d <= 8'hC0; 15'h34FE: d <= 8'hC0; 15'h34FF: d <= 8'hC0;
                15'h3500: d <= 8'hC0; 15'h3501: d <= 8'hC0; 15'h3502: d <= 8'hC0; 15'h3503: d <= 8'hC0;
                15'h3504: d <= 8'hC0; 15'h3505: d <= 8'hC0; 15'h3506: d <= 8'hC0; 15'h3507: d <= 8'hC0;
                15'h3508: d <= 8'hC0; 15'h3509: d <= 8'hC0; 15'h350A: d <= 8'hC0; 15'h350B: d <= 8'hC0;
                15'h350C: d <= 8'hC0; 15'h350D: d <= 8'hC0; 15'h350E: d <= 8'hC0; 15'h350F: d <= 8'hC0;
                15'h3510: d <= 8'hC0; 15'h3511: d <= 8'hC0; 15'h3512: d <= 8'hC0; 15'h3513: d <= 8'hC0;
                15'h3514: d <= 8'hC0; 15'h3515: d <= 8'hC0; 15'h3516: d <= 8'hC0; 15'h3517: d <= 8'hC0;
                15'h3518: d <= 8'hC0; 15'h3519: d <= 8'hC0; 15'h351A: d <= 8'hC0; 15'h351B: d <= 8'hC0;
                15'h351C: d <= 8'hC0; 15'h351D: d <= 8'hC0; 15'h351E: d <= 8'hC0; 15'h351F: d <= 8'hC0;
                15'h3520: d <= 8'hC0; 15'h3521: d <= 8'hC0; 15'h3522: d <= 8'hC0; 15'h3523: d <= 8'hC0;
                15'h3524: d <= 8'hC0; 15'h3525: d <= 8'hC0; 15'h3526: d <= 8'hC0; 15'h3527: d <= 8'hC0;
                15'h3528: d <= 8'hC0; 15'h3529: d <= 8'hC0; 15'h352A: d <= 8'hC0; 15'h352B: d <= 8'hC0;
                15'h352C: d <= 8'hC0; 15'h352D: d <= 8'hC0; 15'h352E: d <= 8'hC0; 15'h352F: d <= 8'hC0;
                15'h3530: d <= 8'hC0; 15'h3531: d <= 8'hC0; 15'h3532: d <= 8'hC0; 15'h3533: d <= 8'hC0;
                15'h3534: d <= 8'hC0; 15'h3535: d <= 8'hC0; 15'h3536: d <= 8'hC0; 15'h3537: d <= 8'hC0;
                15'h3538: d <= 8'hC0; 15'h3539: d <= 8'hC0; 15'h353A: d <= 8'hC0; 15'h353B: d <= 8'hC0;
                15'h353C: d <= 8'hC0; 15'h353D: d <= 8'hC0; 15'h353E: d <= 8'hC0; 15'h353F: d <= 8'hC0;
                15'h3540: d <= 8'hC0; 15'h3541: d <= 8'hC0; 15'h3542: d <= 8'hC0; 15'h3543: d <= 8'hC0;
                15'h3544: d <= 8'hC0; 15'h3545: d <= 8'hC0; 15'h3546: d <= 8'hC0; 15'h3547: d <= 8'hC0;
                15'h3548: d <= 8'hC0; 15'h3549: d <= 8'hC0; 15'h354A: d <= 8'hC0; 15'h354B: d <= 8'hC0;
                15'h354C: d <= 8'hC0; 15'h354D: d <= 8'hC0; 15'h354E: d <= 8'hC0; 15'h354F: d <= 8'hC0;
                15'h3550: d <= 8'hC0; 15'h3551: d <= 8'hC0; 15'h3552: d <= 8'hC0; 15'h3553: d <= 8'hC0;
                15'h3554: d <= 8'hC0; 15'h3555: d <= 8'hC0; 15'h3556: d <= 8'hC0; 15'h3557: d <= 8'hC0;
                15'h3558: d <= 8'hC0; 15'h3559: d <= 8'hC0; 15'h355A: d <= 8'hC0; 15'h355B: d <= 8'hC0;
                15'h355C: d <= 8'hC0; 15'h355D: d <= 8'hC0; 15'h355E: d <= 8'hC0; 15'h355F: d <= 8'hC0;
                15'h3560: d <= 8'hC0; 15'h3561: d <= 8'hC0; 15'h3562: d <= 8'hC0; 15'h3563: d <= 8'hC0;
                15'h3564: d <= 8'hC0; 15'h3565: d <= 8'hC0; 15'h3566: d <= 8'hC0; 15'h3567: d <= 8'hC0;
                15'h3568: d <= 8'hC0; 15'h3569: d <= 8'hC0; 15'h356A: d <= 8'hC0; 15'h356B: d <= 8'hC0;
                15'h356C: d <= 8'hC0; 15'h356D: d <= 8'hC0; 15'h356E: d <= 8'hC0; 15'h356F: d <= 8'hC0;
                15'h3570: d <= 8'hC0; 15'h3571: d <= 8'hC0; 15'h3572: d <= 8'hC0; 15'h3573: d <= 8'hC0;
                15'h3574: d <= 8'hC0; 15'h3575: d <= 8'hC0; 15'h3576: d <= 8'hC0; 15'h3577: d <= 8'hC0;
                15'h3578: d <= 8'hC0; 15'h3579: d <= 8'hC0; 15'h357A: d <= 8'hC0; 15'h357B: d <= 8'hC0;
                15'h357C: d <= 8'hC0; 15'h357D: d <= 8'hC0; 15'h357E: d <= 8'hC0; 15'h357F: d <= 8'hC0;
                15'h3580: d <= 8'hC0; 15'h3581: d <= 8'hC0; 15'h3582: d <= 8'hC0; 15'h3583: d <= 8'hC0;
                15'h3584: d <= 8'hC0; 15'h3585: d <= 8'hC0; 15'h3586: d <= 8'hC0; 15'h3587: d <= 8'hC0;
                15'h3588: d <= 8'hC0; 15'h3589: d <= 8'hC0; 15'h358A: d <= 8'hC0; 15'h358B: d <= 8'hC0;
                15'h358C: d <= 8'hC0; 15'h358D: d <= 8'hC0; 15'h358E: d <= 8'hC0; 15'h358F: d <= 8'hC0;
                15'h3590: d <= 8'hC0; 15'h3591: d <= 8'hC0; 15'h3592: d <= 8'hC0; 15'h3593: d <= 8'hC0;
                15'h3594: d <= 8'hC0; 15'h3595: d <= 8'hC0; 15'h3596: d <= 8'hC0; 15'h3597: d <= 8'hC0;
                15'h3598: d <= 8'hC0; 15'h3599: d <= 8'hC0; 15'h359A: d <= 8'hC0; 15'h359B: d <= 8'hC0;
                15'h359C: d <= 8'hC0; 15'h359D: d <= 8'hC0; 15'h359E: d <= 8'hC0; 15'h359F: d <= 8'hC0;
                15'h35A0: d <= 8'hC0; 15'h35A1: d <= 8'hC0; 15'h35A2: d <= 8'hC0; 15'h35A3: d <= 8'hC0;
                15'h35A4: d <= 8'hC0; 15'h35A5: d <= 8'hC0; 15'h35A6: d <= 8'hC0; 15'h35A7: d <= 8'hC0;
                15'h35A8: d <= 8'hC0; 15'h35A9: d <= 8'hC0; 15'h35AA: d <= 8'hC0; 15'h35AB: d <= 8'hC0;
                15'h35AC: d <= 8'hC0; 15'h35AD: d <= 8'hC0; 15'h35AE: d <= 8'hC0; 15'h35AF: d <= 8'hC0;
                15'h35B0: d <= 8'hC0; 15'h35B1: d <= 8'hC0; 15'h35B2: d <= 8'hC0; 15'h35B3: d <= 8'hC0;
                15'h35B4: d <= 8'hC0; 15'h35B5: d <= 8'hC0; 15'h35B6: d <= 8'hC0; 15'h35B7: d <= 8'hC0;
                15'h35B8: d <= 8'hC0; 15'h35B9: d <= 8'hC0; 15'h35BA: d <= 8'hC0; 15'h35BB: d <= 8'hC0;
                15'h35BC: d <= 8'hC0; 15'h35BD: d <= 8'hC0; 15'h35BE: d <= 8'hC0; 15'h35BF: d <= 8'hC0;
                15'h35C0: d <= 8'hC0; 15'h35C1: d <= 8'hC0; 15'h35C2: d <= 8'hC0; 15'h35C3: d <= 8'hC0;
                15'h35C4: d <= 8'hC0; 15'h35C5: d <= 8'hC0; 15'h35C6: d <= 8'hC0; 15'h35C7: d <= 8'hC0;
                15'h35C8: d <= 8'hC0; 15'h35C9: d <= 8'hC0; 15'h35CA: d <= 8'hC0; 15'h35CB: d <= 8'hC0;
                15'h35CC: d <= 8'hC0; 15'h35CD: d <= 8'hC0; 15'h35CE: d <= 8'hC0; 15'h35CF: d <= 8'hC0;
                15'h35D0: d <= 8'hC0; 15'h35D1: d <= 8'hC0; 15'h35D2: d <= 8'hC0; 15'h35D3: d <= 8'hC0;
                15'h35D4: d <= 8'hC0; 15'h35D5: d <= 8'hC0; 15'h35D6: d <= 8'hC0; 15'h35D7: d <= 8'hC0;
                15'h35D8: d <= 8'hC0; 15'h35D9: d <= 8'hC0; 15'h35DA: d <= 8'hC0; 15'h35DB: d <= 8'hC0;
                15'h35DC: d <= 8'hC0; 15'h35DD: d <= 8'hC0; 15'h35DE: d <= 8'hC0; 15'h35DF: d <= 8'hC0;
                15'h35E0: d <= 8'hC0; 15'h35E1: d <= 8'hC0; 15'h35E2: d <= 8'hC0; 15'h35E3: d <= 8'hC0;
                15'h35E4: d <= 8'hC0; 15'h35E5: d <= 8'hC0; 15'h35E6: d <= 8'hC0; 15'h35E7: d <= 8'hC0;
                15'h35E8: d <= 8'hC0; 15'h35E9: d <= 8'hC0; 15'h35EA: d <= 8'hC0; 15'h35EB: d <= 8'hC0;
                15'h35EC: d <= 8'hC0; 15'h35ED: d <= 8'hC0; 15'h35EE: d <= 8'hC0; 15'h35EF: d <= 8'hC0;
                15'h35F0: d <= 8'hC0; 15'h35F1: d <= 8'hC0; 15'h35F2: d <= 8'hC0; 15'h35F3: d <= 8'hC0;
                15'h35F4: d <= 8'hC0; 15'h35F5: d <= 8'hC0; 15'h35F6: d <= 8'hC0; 15'h35F7: d <= 8'hC0;
                15'h35F8: d <= 8'hC0; 15'h35F9: d <= 8'hC0; 15'h35FA: d <= 8'hC0; 15'h35FB: d <= 8'hC0;
                15'h35FC: d <= 8'hC0; 15'h35FD: d <= 8'hC0; 15'h35FE: d <= 8'hC0; 15'h35FF: d <= 8'hC0;
                15'h3600: d <= 8'hC0; 15'h3601: d <= 8'hC0; 15'h3602: d <= 8'hC0; 15'h3603: d <= 8'hC0;
                15'h3604: d <= 8'hC0; 15'h3605: d <= 8'hC0; 15'h3606: d <= 8'hC0; 15'h3607: d <= 8'hC0;
                15'h3608: d <= 8'hC0; 15'h3609: d <= 8'hC0; 15'h360A: d <= 8'hC0; 15'h360B: d <= 8'hC0;
                15'h360C: d <= 8'hC0; 15'h360D: d <= 8'hC0; 15'h360E: d <= 8'hC0; 15'h360F: d <= 8'hC0;
                15'h3610: d <= 8'hC0; 15'h3611: d <= 8'hC0; 15'h3612: d <= 8'hC0; 15'h3613: d <= 8'hC0;
                15'h3614: d <= 8'hC0; 15'h3615: d <= 8'hC0; 15'h3616: d <= 8'hC0; 15'h3617: d <= 8'hC0;
                15'h3618: d <= 8'hC0; 15'h3619: d <= 8'hC0; 15'h361A: d <= 8'hC0; 15'h361B: d <= 8'hC0;
                15'h361C: d <= 8'hC0; 15'h361D: d <= 8'hC0; 15'h361E: d <= 8'hC0; 15'h361F: d <= 8'hC0;
                15'h3620: d <= 8'hC0; 15'h3621: d <= 8'hC0; 15'h3622: d <= 8'hC0; 15'h3623: d <= 8'hC0;
                15'h3624: d <= 8'hC0; 15'h3625: d <= 8'hC0; 15'h3626: d <= 8'hC0; 15'h3627: d <= 8'hC0;
                15'h3628: d <= 8'hC0; 15'h3629: d <= 8'hC0; 15'h362A: d <= 8'hC0; 15'h362B: d <= 8'hC0;
                15'h362C: d <= 8'hC0; 15'h362D: d <= 8'hC0; 15'h362E: d <= 8'hC0; 15'h362F: d <= 8'hC0;
                15'h3630: d <= 8'hC0; 15'h3631: d <= 8'hC0; 15'h3632: d <= 8'hC0; 15'h3633: d <= 8'hC0;
                15'h3634: d <= 8'hC0; 15'h3635: d <= 8'hC0; 15'h3636: d <= 8'hC0; 15'h3637: d <= 8'hC0;
                15'h3638: d <= 8'hC0; 15'h3639: d <= 8'hC0; 15'h363A: d <= 8'hC0; 15'h363B: d <= 8'hC0;
                15'h363C: d <= 8'hC0; 15'h363D: d <= 8'hC0; 15'h363E: d <= 8'hC0; 15'h363F: d <= 8'hC0;
                15'h3640: d <= 8'hC0; 15'h3641: d <= 8'hC0; 15'h3642: d <= 8'hC0; 15'h3643: d <= 8'hC0;
                15'h3644: d <= 8'hC0; 15'h3645: d <= 8'hC0; 15'h3646: d <= 8'hC0; 15'h3647: d <= 8'hC0;
                15'h3648: d <= 8'hC0; 15'h3649: d <= 8'hC0; 15'h364A: d <= 8'hC0; 15'h364B: d <= 8'hC0;
                15'h364C: d <= 8'hC0; 15'h364D: d <= 8'hC0; 15'h364E: d <= 8'hC0; 15'h364F: d <= 8'hC0;
                15'h3650: d <= 8'hC0; 15'h3651: d <= 8'hC0; 15'h3652: d <= 8'hC0; 15'h3653: d <= 8'hC0;
                15'h3654: d <= 8'hC0; 15'h3655: d <= 8'hC0; 15'h3656: d <= 8'hC0; 15'h3657: d <= 8'hC0;
                15'h3658: d <= 8'hC0; 15'h3659: d <= 8'hC0; 15'h365A: d <= 8'hC0; 15'h365B: d <= 8'hC0;
                15'h365C: d <= 8'hC0; 15'h365D: d <= 8'hC0; 15'h365E: d <= 8'hC0; 15'h365F: d <= 8'hC0;
                15'h3660: d <= 8'hC0; 15'h3661: d <= 8'hC0; 15'h3662: d <= 8'hC0; 15'h3663: d <= 8'hC0;
                15'h3664: d <= 8'hC0; 15'h3665: d <= 8'hC0; 15'h3666: d <= 8'hC0; 15'h3667: d <= 8'hC0;
                15'h3668: d <= 8'hC0; 15'h3669: d <= 8'hC0; 15'h366A: d <= 8'hC0; 15'h366B: d <= 8'hC0;
                15'h366C: d <= 8'hC0; 15'h366D: d <= 8'hC0; 15'h366E: d <= 8'hC0; 15'h366F: d <= 8'hC0;
                15'h3670: d <= 8'hC0; 15'h3671: d <= 8'hC0; 15'h3672: d <= 8'hC0; 15'h3673: d <= 8'hC0;
                15'h3674: d <= 8'hC0; 15'h3675: d <= 8'hC0; 15'h3676: d <= 8'hC0; 15'h3677: d <= 8'hC0;
                15'h3678: d <= 8'hC0; 15'h3679: d <= 8'hC0; 15'h367A: d <= 8'hC0; 15'h367B: d <= 8'hC0;
                15'h367C: d <= 8'hC0; 15'h367D: d <= 8'hC0; 15'h367E: d <= 8'hC0; 15'h367F: d <= 8'hC0;
                15'h3680: d <= 8'hC0; 15'h3681: d <= 8'hC0; 15'h3682: d <= 8'hC0; 15'h3683: d <= 8'hC0;
                15'h3684: d <= 8'hC0; 15'h3685: d <= 8'hC0; 15'h3686: d <= 8'hC0; 15'h3687: d <= 8'hC0;
                15'h3688: d <= 8'hC0; 15'h3689: d <= 8'hC0; 15'h368A: d <= 8'hC0; 15'h368B: d <= 8'hC0;
                15'h368C: d <= 8'hC0; 15'h368D: d <= 8'hC0; 15'h368E: d <= 8'hC0; 15'h368F: d <= 8'hC0;
                15'h3690: d <= 8'hC0; 15'h3691: d <= 8'hC0; 15'h3692: d <= 8'hC0; 15'h3693: d <= 8'hC0;
                15'h3694: d <= 8'hC0; 15'h3695: d <= 8'hC0; 15'h3696: d <= 8'hC0; 15'h3697: d <= 8'hC0;
                15'h3698: d <= 8'hC0; 15'h3699: d <= 8'hC0; 15'h369A: d <= 8'hC0; 15'h369B: d <= 8'hC0;
                15'h369C: d <= 8'hC0; 15'h369D: d <= 8'hC0; 15'h369E: d <= 8'hC0; 15'h369F: d <= 8'hC0;
                15'h36A0: d <= 8'hC0; 15'h36A1: d <= 8'hC0; 15'h36A2: d <= 8'hC0; 15'h36A3: d <= 8'hC0;
                15'h36A4: d <= 8'hC0; 15'h36A5: d <= 8'hC0; 15'h36A6: d <= 8'hC0; 15'h36A7: d <= 8'hC0;
                15'h36A8: d <= 8'hC0; 15'h36A9: d <= 8'hC0; 15'h36AA: d <= 8'hC0; 15'h36AB: d <= 8'hC0;
                15'h36AC: d <= 8'hC0; 15'h36AD: d <= 8'hC0; 15'h36AE: d <= 8'hC0; 15'h36AF: d <= 8'hC0;
                15'h36B0: d <= 8'hC0; 15'h36B1: d <= 8'hC0; 15'h36B2: d <= 8'hC0; 15'h36B3: d <= 8'hC0;
                15'h36B4: d <= 8'hC0; 15'h36B5: d <= 8'hC0; 15'h36B6: d <= 8'hC0; 15'h36B7: d <= 8'hC0;
                15'h36B8: d <= 8'hC0; 15'h36B9: d <= 8'hC0; 15'h36BA: d <= 8'hC0; 15'h36BB: d <= 8'hC0;
                15'h36BC: d <= 8'hC0; 15'h36BD: d <= 8'hC0; 15'h36BE: d <= 8'hC0; 15'h36BF: d <= 8'hC0;
                15'h36C0: d <= 8'hC0; 15'h36C1: d <= 8'hC0; 15'h36C2: d <= 8'hC0; 15'h36C3: d <= 8'hC0;
                15'h36C4: d <= 8'hC0; 15'h36C5: d <= 8'hC0; 15'h36C6: d <= 8'hC0; 15'h36C7: d <= 8'hC0;
                15'h36C8: d <= 8'hC0; 15'h36C9: d <= 8'hC0; 15'h36CA: d <= 8'hC0; 15'h36CB: d <= 8'hC0;
                15'h36CC: d <= 8'hC0; 15'h36CD: d <= 8'hC0; 15'h36CE: d <= 8'hC0; 15'h36CF: d <= 8'hC0;
                15'h36D0: d <= 8'hC0; 15'h36D1: d <= 8'hC0; 15'h36D2: d <= 8'hC0; 15'h36D3: d <= 8'hC0;
                15'h36D4: d <= 8'hC0; 15'h36D5: d <= 8'hC0; 15'h36D6: d <= 8'hC0; 15'h36D7: d <= 8'hC0;
                15'h36D8: d <= 8'hC0; 15'h36D9: d <= 8'hC0; 15'h36DA: d <= 8'hC0; 15'h36DB: d <= 8'hC0;
                15'h36DC: d <= 8'hC0; 15'h36DD: d <= 8'hC0; 15'h36DE: d <= 8'hC0; 15'h36DF: d <= 8'hC0;
                15'h36E0: d <= 8'hC0; 15'h36E1: d <= 8'hC0; 15'h36E2: d <= 8'hC0; 15'h36E3: d <= 8'hC0;
                15'h36E4: d <= 8'hC0; 15'h36E5: d <= 8'hC0; 15'h36E6: d <= 8'hC0; 15'h36E7: d <= 8'hC0;
                15'h36E8: d <= 8'hC0; 15'h36E9: d <= 8'hC0; 15'h36EA: d <= 8'hC0; 15'h36EB: d <= 8'hC0;
                15'h36EC: d <= 8'hC0; 15'h36ED: d <= 8'hC0; 15'h36EE: d <= 8'hC0; 15'h36EF: d <= 8'hC0;
                15'h36F0: d <= 8'hC0; 15'h36F1: d <= 8'hC0; 15'h36F2: d <= 8'hC0; 15'h36F3: d <= 8'hC0;
                15'h36F4: d <= 8'hC0; 15'h36F5: d <= 8'hC0; 15'h36F6: d <= 8'hC0; 15'h36F7: d <= 8'hC0;
                15'h36F8: d <= 8'hC0; 15'h36F9: d <= 8'hC0; 15'h36FA: d <= 8'hC0; 15'h36FB: d <= 8'hC0;
                15'h36FC: d <= 8'hC0; 15'h36FD: d <= 8'hC0; 15'h36FE: d <= 8'hC0; 15'h36FF: d <= 8'hC0;
                15'h3700: d <= 8'hC0; 15'h3701: d <= 8'hC0; 15'h3702: d <= 8'hC0; 15'h3703: d <= 8'hC0;
                15'h3704: d <= 8'hC0; 15'h3705: d <= 8'hC0; 15'h3706: d <= 8'hC0; 15'h3707: d <= 8'hC0;
                15'h3708: d <= 8'hC0; 15'h3709: d <= 8'hC0; 15'h370A: d <= 8'hC0; 15'h370B: d <= 8'hC0;
                15'h370C: d <= 8'hC0; 15'h370D: d <= 8'hC0; 15'h370E: d <= 8'hC0; 15'h370F: d <= 8'hC0;
                15'h3710: d <= 8'hC0; 15'h3711: d <= 8'hC0; 15'h3712: d <= 8'hC0; 15'h3713: d <= 8'hC0;
                15'h3714: d <= 8'hC0; 15'h3715: d <= 8'hC0; 15'h3716: d <= 8'hC0; 15'h3717: d <= 8'hC0;
                15'h3718: d <= 8'hC0; 15'h3719: d <= 8'hC0; 15'h371A: d <= 8'hC0; 15'h371B: d <= 8'hC0;
                15'h371C: d <= 8'hC0; 15'h371D: d <= 8'hC0; 15'h371E: d <= 8'hC0; 15'h371F: d <= 8'hC0;
                15'h3720: d <= 8'hC0; 15'h3721: d <= 8'hC0; 15'h3722: d <= 8'hC0; 15'h3723: d <= 8'hC0;
                15'h3724: d <= 8'hC0; 15'h3725: d <= 8'hC0; 15'h3726: d <= 8'hC0; 15'h3727: d <= 8'hC0;
                15'h3728: d <= 8'hC0; 15'h3729: d <= 8'hC0; 15'h372A: d <= 8'hC0; 15'h372B: d <= 8'hC0;
                15'h372C: d <= 8'hC0; 15'h372D: d <= 8'hC0; 15'h372E: d <= 8'hC0; 15'h372F: d <= 8'hC0;
                15'h3730: d <= 8'hC0; 15'h3731: d <= 8'hC0; 15'h3732: d <= 8'hC0; 15'h3733: d <= 8'hC0;
                15'h3734: d <= 8'hC0; 15'h3735: d <= 8'hC0; 15'h3736: d <= 8'hC0; 15'h3737: d <= 8'hC0;
                15'h3738: d <= 8'hC0; 15'h3739: d <= 8'hC0; 15'h373A: d <= 8'hC0; 15'h373B: d <= 8'hC0;
                15'h373C: d <= 8'hC0; 15'h373D: d <= 8'hC0; 15'h373E: d <= 8'hC0; 15'h373F: d <= 8'hC0;
                15'h3740: d <= 8'hC0; 15'h3741: d <= 8'hC0; 15'h3742: d <= 8'hC0; 15'h3743: d <= 8'hC0;
                15'h3744: d <= 8'hC0; 15'h3745: d <= 8'hC0; 15'h3746: d <= 8'hC0; 15'h3747: d <= 8'hC0;
                15'h3748: d <= 8'hC0; 15'h3749: d <= 8'hC0; 15'h374A: d <= 8'hC0; 15'h374B: d <= 8'hC0;
                15'h374C: d <= 8'hC0; 15'h374D: d <= 8'hC0; 15'h374E: d <= 8'hC0; 15'h374F: d <= 8'hC0;
                15'h3750: d <= 8'hC0; 15'h3751: d <= 8'hC0; 15'h3752: d <= 8'hC0; 15'h3753: d <= 8'hC0;
                15'h3754: d <= 8'hC0; 15'h3755: d <= 8'hC0; 15'h3756: d <= 8'hC0; 15'h3757: d <= 8'hC0;
                15'h3758: d <= 8'hC0; 15'h3759: d <= 8'hC0; 15'h375A: d <= 8'hC0; 15'h375B: d <= 8'hC0;
                15'h375C: d <= 8'hC0; 15'h375D: d <= 8'hC0; 15'h375E: d <= 8'hC0; 15'h375F: d <= 8'hC0;
                15'h3760: d <= 8'hC0; 15'h3761: d <= 8'hC0; 15'h3762: d <= 8'hC0; 15'h3763: d <= 8'hC0;
                15'h3764: d <= 8'hC0; 15'h3765: d <= 8'hC0; 15'h3766: d <= 8'hC0; 15'h3767: d <= 8'hC0;
                15'h3768: d <= 8'hC0; 15'h3769: d <= 8'hC0; 15'h376A: d <= 8'hC0; 15'h376B: d <= 8'hC0;
                15'h376C: d <= 8'hC0; 15'h376D: d <= 8'hC0; 15'h376E: d <= 8'hC0; 15'h376F: d <= 8'hC0;
                15'h3770: d <= 8'hC0; 15'h3771: d <= 8'hC0; 15'h3772: d <= 8'hC0; 15'h3773: d <= 8'hC0;
                15'h3774: d <= 8'hC0; 15'h3775: d <= 8'hC0; 15'h3776: d <= 8'hC0; 15'h3777: d <= 8'hC0;
                15'h3778: d <= 8'hC0; 15'h3779: d <= 8'hC0; 15'h377A: d <= 8'hC0; 15'h377B: d <= 8'hC0;
                15'h377C: d <= 8'hC0; 15'h377D: d <= 8'hC0; 15'h377E: d <= 8'hC0; 15'h377F: d <= 8'hC0;
                15'h3780: d <= 8'hC0; 15'h3781: d <= 8'hC0; 15'h3782: d <= 8'hC0; 15'h3783: d <= 8'hC0;
                15'h3784: d <= 8'hC0; 15'h3785: d <= 8'hC0; 15'h3786: d <= 8'hC0; 15'h3787: d <= 8'hC0;
                15'h3788: d <= 8'hC0; 15'h3789: d <= 8'hC0; 15'h378A: d <= 8'hC0; 15'h378B: d <= 8'hC0;
                15'h378C: d <= 8'hC0; 15'h378D: d <= 8'hC0; 15'h378E: d <= 8'hC0; 15'h378F: d <= 8'hC0;
                15'h3790: d <= 8'hC0; 15'h3791: d <= 8'hC0; 15'h3792: d <= 8'hC0; 15'h3793: d <= 8'hC0;
                15'h3794: d <= 8'hC0; 15'h3795: d <= 8'hC0; 15'h3796: d <= 8'hC0; 15'h3797: d <= 8'hC0;
                15'h3798: d <= 8'hC0; 15'h3799: d <= 8'hC0; 15'h379A: d <= 8'hC0; 15'h379B: d <= 8'hC0;
                15'h379C: d <= 8'hC0; 15'h379D: d <= 8'hC0; 15'h379E: d <= 8'hC0; 15'h379F: d <= 8'hC0;
                15'h37A0: d <= 8'hC0; 15'h37A1: d <= 8'hC0; 15'h37A2: d <= 8'hC0; 15'h37A3: d <= 8'hC0;
                15'h37A4: d <= 8'hC0; 15'h37A5: d <= 8'hC0; 15'h37A6: d <= 8'hC0; 15'h37A7: d <= 8'hC0;
                15'h37A8: d <= 8'hC0; 15'h37A9: d <= 8'hC0; 15'h37AA: d <= 8'hC0; 15'h37AB: d <= 8'hC0;
                15'h37AC: d <= 8'hC0; 15'h37AD: d <= 8'hC0; 15'h37AE: d <= 8'hC0; 15'h37AF: d <= 8'hC0;
                15'h37B0: d <= 8'hC0; 15'h37B1: d <= 8'hC0; 15'h37B2: d <= 8'hC0; 15'h37B3: d <= 8'hC0;
                15'h37B4: d <= 8'hC0; 15'h37B5: d <= 8'hC0; 15'h37B6: d <= 8'hC0; 15'h37B7: d <= 8'hC0;
                15'h37B8: d <= 8'hC0; 15'h37B9: d <= 8'hC0; 15'h37BA: d <= 8'hC0; 15'h37BB: d <= 8'hC0;
                15'h37BC: d <= 8'hC0; 15'h37BD: d <= 8'hC0; 15'h37BE: d <= 8'hC0; 15'h37BF: d <= 8'hC0;
                15'h37C0: d <= 8'hC0; 15'h37C1: d <= 8'hC0; 15'h37C2: d <= 8'hC0; 15'h37C3: d <= 8'hC0;
                15'h37C4: d <= 8'hC0; 15'h37C5: d <= 8'hC0; 15'h37C6: d <= 8'hC0; 15'h37C7: d <= 8'hC0;
                15'h37C8: d <= 8'hC0; 15'h37C9: d <= 8'hC0; 15'h37CA: d <= 8'hC0; 15'h37CB: d <= 8'hC0;
                15'h37CC: d <= 8'hC0; 15'h37CD: d <= 8'hC0; 15'h37CE: d <= 8'hC0; 15'h37CF: d <= 8'hC0;
                15'h37D0: d <= 8'hC0; 15'h37D1: d <= 8'hC0; 15'h37D2: d <= 8'hC0; 15'h37D3: d <= 8'hC0;
                15'h37D4: d <= 8'hC0; 15'h37D5: d <= 8'hC0; 15'h37D6: d <= 8'hC0; 15'h37D7: d <= 8'hC0;
                15'h37D8: d <= 8'hC0; 15'h37D9: d <= 8'hC0; 15'h37DA: d <= 8'hC0; 15'h37DB: d <= 8'hC0;
                15'h37DC: d <= 8'hC0; 15'h37DD: d <= 8'hC0; 15'h37DE: d <= 8'hC0; 15'h37DF: d <= 8'hC0;
                15'h37E0: d <= 8'hC0; 15'h37E1: d <= 8'hC0; 15'h37E2: d <= 8'hC0; 15'h37E3: d <= 8'hC0;
                15'h37E4: d <= 8'hC0; 15'h37E5: d <= 8'hC0; 15'h37E6: d <= 8'hC0; 15'h37E7: d <= 8'hC0;
                15'h37E8: d <= 8'hC0; 15'h37E9: d <= 8'hC0; 15'h37EA: d <= 8'hC0; 15'h37EB: d <= 8'hC0;
                15'h37EC: d <= 8'hC0; 15'h37ED: d <= 8'hC0; 15'h37EE: d <= 8'hC0; 15'h37EF: d <= 8'hC0;
                15'h37F0: d <= 8'hC0; 15'h37F1: d <= 8'hC0; 15'h37F2: d <= 8'hC0; 15'h37F3: d <= 8'hC0;
                15'h37F4: d <= 8'hC0; 15'h37F5: d <= 8'hC0; 15'h37F6: d <= 8'hC0; 15'h37F7: d <= 8'hC0;
                15'h37F8: d <= 8'hC0; 15'h37F9: d <= 8'hC0; 15'h37FA: d <= 8'hC0; 15'h37FB: d <= 8'hC0;
                15'h37FC: d <= 8'hC0; 15'h37FD: d <= 8'hC0; 15'h37FE: d <= 8'hC0; 15'h37FF: d <= 8'hC0;
                15'h3800: d <= 8'hC0; 15'h3801: d <= 8'hC0; 15'h3802: d <= 8'hC0; 15'h3803: d <= 8'hC0;
                15'h3804: d <= 8'hC0; 15'h3805: d <= 8'hC0; 15'h3806: d <= 8'hC0; 15'h3807: d <= 8'hC0;
                15'h3808: d <= 8'hC0; 15'h3809: d <= 8'hC0; 15'h380A: d <= 8'hC0; 15'h380B: d <= 8'hC0;
                15'h380C: d <= 8'hC0; 15'h380D: d <= 8'hC0; 15'h380E: d <= 8'hC0; 15'h380F: d <= 8'hC0;
                15'h3810: d <= 8'hC0; 15'h3811: d <= 8'hC0; 15'h3812: d <= 8'hC0; 15'h3813: d <= 8'hC0;
                15'h3814: d <= 8'hC0; 15'h3815: d <= 8'hC0; 15'h3816: d <= 8'hC0; 15'h3817: d <= 8'hC0;
                15'h3818: d <= 8'hC0; 15'h3819: d <= 8'hC0; 15'h381A: d <= 8'hC0; 15'h381B: d <= 8'hC0;
                15'h381C: d <= 8'hC0; 15'h381D: d <= 8'hC0; 15'h381E: d <= 8'hC0; 15'h381F: d <= 8'hC0;
                15'h3820: d <= 8'hC0; 15'h3821: d <= 8'hC0; 15'h3822: d <= 8'hC0; 15'h3823: d <= 8'hC0;
                15'h3824: d <= 8'hC0; 15'h3825: d <= 8'hC0; 15'h3826: d <= 8'hC0; 15'h3827: d <= 8'hC0;
                15'h3828: d <= 8'hC0; 15'h3829: d <= 8'hC0; 15'h382A: d <= 8'hC0; 15'h382B: d <= 8'hC0;
                15'h382C: d <= 8'hC0; 15'h382D: d <= 8'hC0; 15'h382E: d <= 8'hC0; 15'h382F: d <= 8'hC0;
                15'h3830: d <= 8'hC0; 15'h3831: d <= 8'hC0; 15'h3832: d <= 8'hC0; 15'h3833: d <= 8'hC0;
                15'h3834: d <= 8'hC0; 15'h3835: d <= 8'hC0; 15'h3836: d <= 8'hC0; 15'h3837: d <= 8'hC0;
                15'h3838: d <= 8'hC0; 15'h3839: d <= 8'hC0; 15'h383A: d <= 8'hC0; 15'h383B: d <= 8'hC0;
                15'h383C: d <= 8'hC0; 15'h383D: d <= 8'hC0; 15'h383E: d <= 8'hC0; 15'h383F: d <= 8'hC0;
                15'h3840: d <= 8'hC0; 15'h3841: d <= 8'hC0; 15'h3842: d <= 8'hC0; 15'h3843: d <= 8'hC0;
                15'h3844: d <= 8'hC0; 15'h3845: d <= 8'hC0; 15'h3846: d <= 8'hC0; 15'h3847: d <= 8'hC0;
                15'h3848: d <= 8'hC0; 15'h3849: d <= 8'hC0; 15'h384A: d <= 8'hC0; 15'h384B: d <= 8'hC0;
                15'h384C: d <= 8'hC0; 15'h384D: d <= 8'hC0; 15'h384E: d <= 8'hC0; 15'h384F: d <= 8'hC0;
                15'h3850: d <= 8'hC0; 15'h3851: d <= 8'hC0; 15'h3852: d <= 8'hC0; 15'h3853: d <= 8'hC0;
                15'h3854: d <= 8'hC0; 15'h3855: d <= 8'hC0; 15'h3856: d <= 8'hC0; 15'h3857: d <= 8'hC0;
                15'h3858: d <= 8'hC0; 15'h3859: d <= 8'hC0; 15'h385A: d <= 8'hC0; 15'h385B: d <= 8'hC0;
                15'h385C: d <= 8'hC0; 15'h385D: d <= 8'hC0; 15'h385E: d <= 8'hC0; 15'h385F: d <= 8'hC0;
                15'h3860: d <= 8'hC0; 15'h3861: d <= 8'hC0; 15'h3862: d <= 8'hC0; 15'h3863: d <= 8'hC0;
                15'h3864: d <= 8'hC0; 15'h3865: d <= 8'hC0; 15'h3866: d <= 8'hC0; 15'h3867: d <= 8'hC0;
                15'h3868: d <= 8'hC0; 15'h3869: d <= 8'hC0; 15'h386A: d <= 8'hC0; 15'h386B: d <= 8'hC0;
                15'h386C: d <= 8'hC0; 15'h386D: d <= 8'hC0; 15'h386E: d <= 8'hC0; 15'h386F: d <= 8'hC0;
                15'h3870: d <= 8'hC0; 15'h3871: d <= 8'hC0; 15'h3872: d <= 8'hC0; 15'h3873: d <= 8'hC0;
                15'h3874: d <= 8'hC0; 15'h3875: d <= 8'hC0; 15'h3876: d <= 8'hC0; 15'h3877: d <= 8'hC0;
                15'h3878: d <= 8'hC0; 15'h3879: d <= 8'hC0; 15'h387A: d <= 8'hC0; 15'h387B: d <= 8'hC0;
                15'h387C: d <= 8'hC0; 15'h387D: d <= 8'hC0; 15'h387E: d <= 8'hC0; 15'h387F: d <= 8'hC0;
                15'h3880: d <= 8'hC0; 15'h3881: d <= 8'hC0; 15'h3882: d <= 8'hC0; 15'h3883: d <= 8'hC0;
                15'h3884: d <= 8'hC0; 15'h3885: d <= 8'hC0; 15'h3886: d <= 8'hC0; 15'h3887: d <= 8'hC0;
                15'h3888: d <= 8'hC0; 15'h3889: d <= 8'hC0; 15'h388A: d <= 8'hC0; 15'h388B: d <= 8'hC0;
                15'h388C: d <= 8'hC0; 15'h388D: d <= 8'hC0; 15'h388E: d <= 8'hC0; 15'h388F: d <= 8'hC0;
                15'h3890: d <= 8'hC0; 15'h3891: d <= 8'hC0; 15'h3892: d <= 8'hC0; 15'h3893: d <= 8'hC0;
                15'h3894: d <= 8'hC0; 15'h3895: d <= 8'hC0; 15'h3896: d <= 8'hC0; 15'h3897: d <= 8'hC0;
                15'h3898: d <= 8'hC0; 15'h3899: d <= 8'hC0; 15'h389A: d <= 8'hC0; 15'h389B: d <= 8'hC0;
                15'h389C: d <= 8'hC0; 15'h389D: d <= 8'hC0; 15'h389E: d <= 8'hC0; 15'h389F: d <= 8'hC0;
                15'h38A0: d <= 8'hC0; 15'h38A1: d <= 8'hC0; 15'h38A2: d <= 8'hC0; 15'h38A3: d <= 8'hC0;
                15'h38A4: d <= 8'hC0; 15'h38A5: d <= 8'hC0; 15'h38A6: d <= 8'hC0; 15'h38A7: d <= 8'hC0;
                15'h38A8: d <= 8'hC0; 15'h38A9: d <= 8'hC0; 15'h38AA: d <= 8'hC0; 15'h38AB: d <= 8'hC0;
                15'h38AC: d <= 8'hC0; 15'h38AD: d <= 8'hC0; 15'h38AE: d <= 8'hC0; 15'h38AF: d <= 8'hC0;
                15'h38B0: d <= 8'hC0; 15'h38B1: d <= 8'hC0; 15'h38B2: d <= 8'hC0; 15'h38B3: d <= 8'hC0;
                15'h38B4: d <= 8'hC0; 15'h38B5: d <= 8'hC0; 15'h38B6: d <= 8'hC0; 15'h38B7: d <= 8'hC0;
                15'h38B8: d <= 8'hC0; 15'h38B9: d <= 8'hC0; 15'h38BA: d <= 8'hC0; 15'h38BB: d <= 8'hC0;
                15'h38BC: d <= 8'hC0; 15'h38BD: d <= 8'hC0; 15'h38BE: d <= 8'hC0; 15'h38BF: d <= 8'hC0;
                15'h38C0: d <= 8'hC0; 15'h38C1: d <= 8'hC0; 15'h38C2: d <= 8'hC0; 15'h38C3: d <= 8'hC0;
                15'h38C4: d <= 8'hC0; 15'h38C5: d <= 8'hC0; 15'h38C6: d <= 8'hC0; 15'h38C7: d <= 8'hC0;
                15'h38C8: d <= 8'hC0; 15'h38C9: d <= 8'hC0; 15'h38CA: d <= 8'hC0; 15'h38CB: d <= 8'hC0;
                15'h38CC: d <= 8'hC0; 15'h38CD: d <= 8'hC0; 15'h38CE: d <= 8'hC0; 15'h38CF: d <= 8'hC0;
                15'h38D0: d <= 8'hC0; 15'h38D1: d <= 8'hC0; 15'h38D2: d <= 8'hC0; 15'h38D3: d <= 8'hC0;
                15'h38D4: d <= 8'hC0; 15'h38D5: d <= 8'hC0; 15'h38D6: d <= 8'hC0; 15'h38D7: d <= 8'hC0;
                15'h38D8: d <= 8'hC0; 15'h38D9: d <= 8'hC0; 15'h38DA: d <= 8'hC0; 15'h38DB: d <= 8'hC0;
                15'h38DC: d <= 8'hC0; 15'h38DD: d <= 8'hC0; 15'h38DE: d <= 8'hC0; 15'h38DF: d <= 8'hC0;
                15'h38E0: d <= 8'hC0; 15'h38E1: d <= 8'hC0; 15'h38E2: d <= 8'hC0; 15'h38E3: d <= 8'hC0;
                15'h38E4: d <= 8'hC0; 15'h38E5: d <= 8'hC0; 15'h38E6: d <= 8'hC0; 15'h38E7: d <= 8'hC0;
                15'h38E8: d <= 8'hC0; 15'h38E9: d <= 8'hC0; 15'h38EA: d <= 8'hC0; 15'h38EB: d <= 8'hC0;
                15'h38EC: d <= 8'hC0; 15'h38ED: d <= 8'hC0; 15'h38EE: d <= 8'hC0; 15'h38EF: d <= 8'hC0;
                15'h38F0: d <= 8'hC0; 15'h38F1: d <= 8'hC0; 15'h38F2: d <= 8'hC0; 15'h38F3: d <= 8'hC0;
                15'h38F4: d <= 8'hC0; 15'h38F5: d <= 8'hC0; 15'h38F6: d <= 8'hC0; 15'h38F7: d <= 8'hC0;
                15'h38F8: d <= 8'hC0; 15'h38F9: d <= 8'hC0; 15'h38FA: d <= 8'hC0; 15'h38FB: d <= 8'hC0;
                15'h38FC: d <= 8'hC0; 15'h38FD: d <= 8'hC0; 15'h38FE: d <= 8'hC0; 15'h38FF: d <= 8'hC0;
                15'h3900: d <= 8'hC0; 15'h3901: d <= 8'hC0; 15'h3902: d <= 8'hC0; 15'h3903: d <= 8'hC0;
                15'h3904: d <= 8'hC0; 15'h3905: d <= 8'hC0; 15'h3906: d <= 8'hC0; 15'h3907: d <= 8'hC0;
                15'h3908: d <= 8'hC0; 15'h3909: d <= 8'hC0; 15'h390A: d <= 8'hC0; 15'h390B: d <= 8'hC0;
                15'h390C: d <= 8'hC0; 15'h390D: d <= 8'hC0; 15'h390E: d <= 8'hC0; 15'h390F: d <= 8'hC0;
                15'h3910: d <= 8'hC0; 15'h3911: d <= 8'hC0; 15'h3912: d <= 8'hC0; 15'h3913: d <= 8'hC0;
                15'h3914: d <= 8'hC0; 15'h3915: d <= 8'hC0; 15'h3916: d <= 8'hC0; 15'h3917: d <= 8'hC0;
                15'h3918: d <= 8'hC0; 15'h3919: d <= 8'hC0; 15'h391A: d <= 8'hC0; 15'h391B: d <= 8'hC0;
                15'h391C: d <= 8'hC0; 15'h391D: d <= 8'hC0; 15'h391E: d <= 8'hC0; 15'h391F: d <= 8'hC0;
                15'h3920: d <= 8'hC0; 15'h3921: d <= 8'hC0; 15'h3922: d <= 8'hC0; 15'h3923: d <= 8'hC0;
                15'h3924: d <= 8'hC0; 15'h3925: d <= 8'hC0; 15'h3926: d <= 8'hC0; 15'h3927: d <= 8'hC0;
                15'h3928: d <= 8'hC0; 15'h3929: d <= 8'hC0; 15'h392A: d <= 8'hC0; 15'h392B: d <= 8'hC0;
                15'h392C: d <= 8'hC0; 15'h392D: d <= 8'hC0; 15'h392E: d <= 8'hC0; 15'h392F: d <= 8'hC0;
                15'h3930: d <= 8'hC0; 15'h3931: d <= 8'hC0; 15'h3932: d <= 8'hC0; 15'h3933: d <= 8'hC0;
                15'h3934: d <= 8'hC0; 15'h3935: d <= 8'hC0; 15'h3936: d <= 8'hC0; 15'h3937: d <= 8'hC0;
                15'h3938: d <= 8'hC0; 15'h3939: d <= 8'hC0; 15'h393A: d <= 8'hC0; 15'h393B: d <= 8'hC0;
                15'h393C: d <= 8'hC0; 15'h393D: d <= 8'hC0; 15'h393E: d <= 8'hC0; 15'h393F: d <= 8'hC0;
                15'h3940: d <= 8'hC0; 15'h3941: d <= 8'hC0; 15'h3942: d <= 8'hC0; 15'h3943: d <= 8'hC0;
                15'h3944: d <= 8'hC0; 15'h3945: d <= 8'hC0; 15'h3946: d <= 8'hC0; 15'h3947: d <= 8'hC0;
                15'h3948: d <= 8'hC0; 15'h3949: d <= 8'hC0; 15'h394A: d <= 8'hC0; 15'h394B: d <= 8'hC0;
                15'h394C: d <= 8'hC0; 15'h394D: d <= 8'hC0; 15'h394E: d <= 8'hC0; 15'h394F: d <= 8'hC0;
                15'h3950: d <= 8'hC0; 15'h3951: d <= 8'hC0; 15'h3952: d <= 8'hC0; 15'h3953: d <= 8'hC0;
                15'h3954: d <= 8'hC0; 15'h3955: d <= 8'hC0; 15'h3956: d <= 8'hC0; 15'h3957: d <= 8'hC0;
                15'h3958: d <= 8'hC0; 15'h3959: d <= 8'hC0; 15'h395A: d <= 8'hC0; 15'h395B: d <= 8'hC0;
                15'h395C: d <= 8'hC0; 15'h395D: d <= 8'hC0; 15'h395E: d <= 8'hC0; 15'h395F: d <= 8'hC0;
                15'h3960: d <= 8'hC0; 15'h3961: d <= 8'hC0; 15'h3962: d <= 8'hC0; 15'h3963: d <= 8'hC0;
                15'h3964: d <= 8'hC0; 15'h3965: d <= 8'hC0; 15'h3966: d <= 8'hC0; 15'h3967: d <= 8'hC0;
                15'h3968: d <= 8'hC0; 15'h3969: d <= 8'hC0; 15'h396A: d <= 8'hC0; 15'h396B: d <= 8'hC0;
                15'h396C: d <= 8'hC0; 15'h396D: d <= 8'hC0; 15'h396E: d <= 8'hC0; 15'h396F: d <= 8'hC0;
                15'h3970: d <= 8'hC0; 15'h3971: d <= 8'hC0; 15'h3972: d <= 8'hC0; 15'h3973: d <= 8'hC0;
                15'h3974: d <= 8'hC0; 15'h3975: d <= 8'hC0; 15'h3976: d <= 8'hC0; 15'h3977: d <= 8'hC0;
                15'h3978: d <= 8'hC0; 15'h3979: d <= 8'hC0; 15'h397A: d <= 8'hC0; 15'h397B: d <= 8'hC0;
                15'h397C: d <= 8'hC0; 15'h397D: d <= 8'hC0; 15'h397E: d <= 8'hC0; 15'h397F: d <= 8'hC0;
                15'h3980: d <= 8'hC0; 15'h3981: d <= 8'hC0; 15'h3982: d <= 8'hC0; 15'h3983: d <= 8'hC0;
                15'h3984: d <= 8'hC0; 15'h3985: d <= 8'hC0; 15'h3986: d <= 8'hC0; 15'h3987: d <= 8'hC0;
                15'h3988: d <= 8'hC0; 15'h3989: d <= 8'hC0; 15'h398A: d <= 8'hC0; 15'h398B: d <= 8'hC0;
                15'h398C: d <= 8'hC0; 15'h398D: d <= 8'hC0; 15'h398E: d <= 8'hC0; 15'h398F: d <= 8'hC0;
                15'h3990: d <= 8'hC0; 15'h3991: d <= 8'hC0; 15'h3992: d <= 8'hC0; 15'h3993: d <= 8'hC0;
                15'h3994: d <= 8'hC0; 15'h3995: d <= 8'hC0; 15'h3996: d <= 8'hC0; 15'h3997: d <= 8'hC0;
                15'h3998: d <= 8'hC0; 15'h3999: d <= 8'hC0; 15'h399A: d <= 8'hC0; 15'h399B: d <= 8'hC0;
                15'h399C: d <= 8'hC0; 15'h399D: d <= 8'hC0; 15'h399E: d <= 8'hC0; 15'h399F: d <= 8'hC0;
                15'h39A0: d <= 8'hC0; 15'h39A1: d <= 8'hC0; 15'h39A2: d <= 8'hC0; 15'h39A3: d <= 8'hC0;
                15'h39A4: d <= 8'hC0; 15'h39A5: d <= 8'hC0; 15'h39A6: d <= 8'hC0; 15'h39A7: d <= 8'hC0;
                15'h39A8: d <= 8'hC0; 15'h39A9: d <= 8'hC0; 15'h39AA: d <= 8'hC0; 15'h39AB: d <= 8'hC0;
                15'h39AC: d <= 8'hC0; 15'h39AD: d <= 8'hC0; 15'h39AE: d <= 8'hC0; 15'h39AF: d <= 8'hC0;
                15'h39B0: d <= 8'hC0; 15'h39B1: d <= 8'hC0; 15'h39B2: d <= 8'hC0; 15'h39B3: d <= 8'hC0;
                15'h39B4: d <= 8'hC0; 15'h39B5: d <= 8'hC0; 15'h39B6: d <= 8'hC0; 15'h39B7: d <= 8'hC0;
                15'h39B8: d <= 8'hC0; 15'h39B9: d <= 8'hC0; 15'h39BA: d <= 8'hC0; 15'h39BB: d <= 8'hC0;
                15'h39BC: d <= 8'hC0; 15'h39BD: d <= 8'hC0; 15'h39BE: d <= 8'hC0; 15'h39BF: d <= 8'hC0;
                15'h39C0: d <= 8'hC0; 15'h39C1: d <= 8'hC0; 15'h39C2: d <= 8'hC0; 15'h39C3: d <= 8'hC0;
                15'h39C4: d <= 8'hC0; 15'h39C5: d <= 8'hC0; 15'h39C6: d <= 8'hC0; 15'h39C7: d <= 8'hC0;
                15'h39C8: d <= 8'hC0; 15'h39C9: d <= 8'hC0; 15'h39CA: d <= 8'hC0; 15'h39CB: d <= 8'hC0;
                15'h39CC: d <= 8'hC0; 15'h39CD: d <= 8'hC0; 15'h39CE: d <= 8'hC0; 15'h39CF: d <= 8'hC0;
                15'h39D0: d <= 8'hC0; 15'h39D1: d <= 8'hC0; 15'h39D2: d <= 8'hC0; 15'h39D3: d <= 8'hC0;
                15'h39D4: d <= 8'hC0; 15'h39D5: d <= 8'hC0; 15'h39D6: d <= 8'hC0; 15'h39D7: d <= 8'hC0;
                15'h39D8: d <= 8'hC0; 15'h39D9: d <= 8'hC0; 15'h39DA: d <= 8'hC0; 15'h39DB: d <= 8'hC0;
                15'h39DC: d <= 8'hC0; 15'h39DD: d <= 8'hC0; 15'h39DE: d <= 8'hC0; 15'h39DF: d <= 8'hC0;
                15'h39E0: d <= 8'hC0; 15'h39E1: d <= 8'hC0; 15'h39E2: d <= 8'hC0; 15'h39E3: d <= 8'hC0;
                15'h39E4: d <= 8'hC0; 15'h39E5: d <= 8'hC0; 15'h39E6: d <= 8'hC0; 15'h39E7: d <= 8'hC0;
                15'h39E8: d <= 8'hC0; 15'h39E9: d <= 8'hC0; 15'h39EA: d <= 8'hC0; 15'h39EB: d <= 8'hC0;
                15'h39EC: d <= 8'hC0; 15'h39ED: d <= 8'hC0; 15'h39EE: d <= 8'hC0; 15'h39EF: d <= 8'hC0;
                15'h39F0: d <= 8'hC0; 15'h39F1: d <= 8'hC0; 15'h39F2: d <= 8'hC0; 15'h39F3: d <= 8'hC0;
                15'h39F4: d <= 8'hC0; 15'h39F5: d <= 8'hC0; 15'h39F6: d <= 8'hC0; 15'h39F7: d <= 8'hC0;
                15'h39F8: d <= 8'hC0; 15'h39F9: d <= 8'hC0; 15'h39FA: d <= 8'hC0; 15'h39FB: d <= 8'hC0;
                15'h39FC: d <= 8'hC0; 15'h39FD: d <= 8'hC0; 15'h39FE: d <= 8'hC0; 15'h39FF: d <= 8'hC0;
                15'h3A00: d <= 8'hC0; 15'h3A01: d <= 8'hC0; 15'h3A02: d <= 8'hC0; 15'h3A03: d <= 8'hC0;
                15'h3A04: d <= 8'hC0; 15'h3A05: d <= 8'hC0; 15'h3A06: d <= 8'hC0; 15'h3A07: d <= 8'hC0;
                15'h3A08: d <= 8'hC0; 15'h3A09: d <= 8'hC0; 15'h3A0A: d <= 8'hC0; 15'h3A0B: d <= 8'hC0;
                15'h3A0C: d <= 8'hC0; 15'h3A0D: d <= 8'hC0; 15'h3A0E: d <= 8'hC0; 15'h3A0F: d <= 8'hC0;
                15'h3A10: d <= 8'hC0; 15'h3A11: d <= 8'hC0; 15'h3A12: d <= 8'hC0; 15'h3A13: d <= 8'hC0;
                15'h3A14: d <= 8'hC0; 15'h3A15: d <= 8'hC0; 15'h3A16: d <= 8'hC0; 15'h3A17: d <= 8'hC0;
                15'h3A18: d <= 8'hC0; 15'h3A19: d <= 8'hC0; 15'h3A1A: d <= 8'hC0; 15'h3A1B: d <= 8'hC0;
                15'h3A1C: d <= 8'hC0; 15'h3A1D: d <= 8'hC0; 15'h3A1E: d <= 8'hC0; 15'h3A1F: d <= 8'hC0;
                15'h3A20: d <= 8'hC0; 15'h3A21: d <= 8'hC0; 15'h3A22: d <= 8'hC0; 15'h3A23: d <= 8'hC0;
                15'h3A24: d <= 8'hC0; 15'h3A25: d <= 8'hC0; 15'h3A26: d <= 8'hC0; 15'h3A27: d <= 8'hC0;
                15'h3A28: d <= 8'hC0; 15'h3A29: d <= 8'hC0; 15'h3A2A: d <= 8'hC0; 15'h3A2B: d <= 8'hC0;
                15'h3A2C: d <= 8'hC0; 15'h3A2D: d <= 8'hC0; 15'h3A2E: d <= 8'hC0; 15'h3A2F: d <= 8'hC0;
                15'h3A30: d <= 8'hC0; 15'h3A31: d <= 8'hC0; 15'h3A32: d <= 8'hC0; 15'h3A33: d <= 8'hC0;
                15'h3A34: d <= 8'hC0; 15'h3A35: d <= 8'hC0; 15'h3A36: d <= 8'hC0; 15'h3A37: d <= 8'hC0;
                15'h3A38: d <= 8'hC0; 15'h3A39: d <= 8'hC0; 15'h3A3A: d <= 8'hC0; 15'h3A3B: d <= 8'hC0;
                15'h3A3C: d <= 8'hC0; 15'h3A3D: d <= 8'hC0; 15'h3A3E: d <= 8'hC0; 15'h3A3F: d <= 8'hC0;
                15'h3A40: d <= 8'hC0; 15'h3A41: d <= 8'hC0; 15'h3A42: d <= 8'hC0; 15'h3A43: d <= 8'hC0;
                15'h3A44: d <= 8'hC0; 15'h3A45: d <= 8'hC0; 15'h3A46: d <= 8'hC0; 15'h3A47: d <= 8'hC0;
                15'h3A48: d <= 8'hC0; 15'h3A49: d <= 8'hC0; 15'h3A4A: d <= 8'hC0; 15'h3A4B: d <= 8'hC0;
                15'h3A4C: d <= 8'hC0; 15'h3A4D: d <= 8'hC0; 15'h3A4E: d <= 8'hC0; 15'h3A4F: d <= 8'hC0;
                15'h3A50: d <= 8'hC0; 15'h3A51: d <= 8'hC0; 15'h3A52: d <= 8'hC0; 15'h3A53: d <= 8'hC0;
                15'h3A54: d <= 8'hC0; 15'h3A55: d <= 8'hC0; 15'h3A56: d <= 8'hC0; 15'h3A57: d <= 8'hC0;
                15'h3A58: d <= 8'hC0; 15'h3A59: d <= 8'hC0; 15'h3A5A: d <= 8'hC0; 15'h3A5B: d <= 8'hC0;
                15'h3A5C: d <= 8'hC0; 15'h3A5D: d <= 8'hC0; 15'h3A5E: d <= 8'hC0; 15'h3A5F: d <= 8'hC0;
                15'h3A60: d <= 8'hC0; 15'h3A61: d <= 8'hC0; 15'h3A62: d <= 8'hC0; 15'h3A63: d <= 8'hC0;
                15'h3A64: d <= 8'hC0; 15'h3A65: d <= 8'hC0; 15'h3A66: d <= 8'hC0; 15'h3A67: d <= 8'hC0;
                15'h3A68: d <= 8'hC0; 15'h3A69: d <= 8'hC0; 15'h3A6A: d <= 8'hC0; 15'h3A6B: d <= 8'hC0;
                15'h3A6C: d <= 8'hC0; 15'h3A6D: d <= 8'hC0; 15'h3A6E: d <= 8'hC0; 15'h3A6F: d <= 8'hC0;
                15'h3A70: d <= 8'hC0; 15'h3A71: d <= 8'hC0; 15'h3A72: d <= 8'hC0; 15'h3A73: d <= 8'hC0;
                15'h3A74: d <= 8'hC0; 15'h3A75: d <= 8'hC0; 15'h3A76: d <= 8'hC0; 15'h3A77: d <= 8'hC0;
                15'h3A78: d <= 8'hC0; 15'h3A79: d <= 8'hC0; 15'h3A7A: d <= 8'hC0; 15'h3A7B: d <= 8'hC0;
                15'h3A7C: d <= 8'hC0; 15'h3A7D: d <= 8'hC0; 15'h3A7E: d <= 8'hC0; 15'h3A7F: d <= 8'hC0;
                15'h3A80: d <= 8'hC0; 15'h3A81: d <= 8'hC0; 15'h3A82: d <= 8'hC0; 15'h3A83: d <= 8'hC0;
                15'h3A84: d <= 8'hC0; 15'h3A85: d <= 8'hC0; 15'h3A86: d <= 8'hC0; 15'h3A87: d <= 8'hC0;
                15'h3A88: d <= 8'hC0; 15'h3A89: d <= 8'hC0; 15'h3A8A: d <= 8'hC0; 15'h3A8B: d <= 8'hC0;
                15'h3A8C: d <= 8'hC0; 15'h3A8D: d <= 8'hC0; 15'h3A8E: d <= 8'hC0; 15'h3A8F: d <= 8'hC0;
                15'h3A90: d <= 8'hC0; 15'h3A91: d <= 8'hC0; 15'h3A92: d <= 8'hC0; 15'h3A93: d <= 8'hC0;
                15'h3A94: d <= 8'hC0; 15'h3A95: d <= 8'hC0; 15'h3A96: d <= 8'hC0; 15'h3A97: d <= 8'hC0;
                15'h3A98: d <= 8'hC0; 15'h3A99: d <= 8'hC0; 15'h3A9A: d <= 8'hC0; 15'h3A9B: d <= 8'hC0;
                15'h3A9C: d <= 8'hC0; 15'h3A9D: d <= 8'hC0; 15'h3A9E: d <= 8'hC0; 15'h3A9F: d <= 8'hC0;
                15'h3AA0: d <= 8'hC0; 15'h3AA1: d <= 8'hC0; 15'h3AA2: d <= 8'hC0; 15'h3AA3: d <= 8'hC0;
                15'h3AA4: d <= 8'hC0; 15'h3AA5: d <= 8'hC0; 15'h3AA6: d <= 8'hC0; 15'h3AA7: d <= 8'hC0;
                15'h3AA8: d <= 8'hC0; 15'h3AA9: d <= 8'hC0; 15'h3AAA: d <= 8'hC0; 15'h3AAB: d <= 8'hC0;
                15'h3AAC: d <= 8'hC0; 15'h3AAD: d <= 8'hC0; 15'h3AAE: d <= 8'hC0; 15'h3AAF: d <= 8'hC0;
                15'h3AB0: d <= 8'hC0; 15'h3AB1: d <= 8'hC0; 15'h3AB2: d <= 8'hC0; 15'h3AB3: d <= 8'hC0;
                15'h3AB4: d <= 8'hC0; 15'h3AB5: d <= 8'hC0; 15'h3AB6: d <= 8'hC0; 15'h3AB7: d <= 8'hC0;
                15'h3AB8: d <= 8'hC0; 15'h3AB9: d <= 8'hC0; 15'h3ABA: d <= 8'hC0; 15'h3ABB: d <= 8'hC0;
                15'h3ABC: d <= 8'hC0; 15'h3ABD: d <= 8'hC0; 15'h3ABE: d <= 8'hC0; 15'h3ABF: d <= 8'hC0;
                15'h3AC0: d <= 8'hC0; 15'h3AC1: d <= 8'hC0; 15'h3AC2: d <= 8'hC0; 15'h3AC3: d <= 8'hC0;
                15'h3AC4: d <= 8'hC0; 15'h3AC5: d <= 8'hC0; 15'h3AC6: d <= 8'hC0; 15'h3AC7: d <= 8'hC0;
                15'h3AC8: d <= 8'hC0; 15'h3AC9: d <= 8'hC0; 15'h3ACA: d <= 8'hC0; 15'h3ACB: d <= 8'hC0;
                15'h3ACC: d <= 8'hC0; 15'h3ACD: d <= 8'hC0; 15'h3ACE: d <= 8'hC0; 15'h3ACF: d <= 8'hC0;
                15'h3AD0: d <= 8'hC0; 15'h3AD1: d <= 8'hC0; 15'h3AD2: d <= 8'hC0; 15'h3AD3: d <= 8'hC0;
                15'h3AD4: d <= 8'hC0; 15'h3AD5: d <= 8'hC0; 15'h3AD6: d <= 8'hC0; 15'h3AD7: d <= 8'hC0;
                15'h3AD8: d <= 8'hC0; 15'h3AD9: d <= 8'hC0; 15'h3ADA: d <= 8'hC0; 15'h3ADB: d <= 8'hC0;
                15'h3ADC: d <= 8'hC0; 15'h3ADD: d <= 8'hC0; 15'h3ADE: d <= 8'hC0; 15'h3ADF: d <= 8'hC0;
                15'h3AE0: d <= 8'hC0; 15'h3AE1: d <= 8'hC0; 15'h3AE2: d <= 8'hC0; 15'h3AE3: d <= 8'hC0;
                15'h3AE4: d <= 8'hC0; 15'h3AE5: d <= 8'hC0; 15'h3AE6: d <= 8'hC0; 15'h3AE7: d <= 8'hC0;
                15'h3AE8: d <= 8'hC0; 15'h3AE9: d <= 8'hC0; 15'h3AEA: d <= 8'hC0; 15'h3AEB: d <= 8'hC0;
                15'h3AEC: d <= 8'hC0; 15'h3AED: d <= 8'hC0; 15'h3AEE: d <= 8'hC0; 15'h3AEF: d <= 8'hC0;
                15'h3AF0: d <= 8'hC0; 15'h3AF1: d <= 8'hC0; 15'h3AF2: d <= 8'hC0; 15'h3AF3: d <= 8'hC0;
                15'h3AF4: d <= 8'hC0; 15'h3AF5: d <= 8'hC0; 15'h3AF6: d <= 8'hC0; 15'h3AF7: d <= 8'hC0;
                15'h3AF8: d <= 8'hC0; 15'h3AF9: d <= 8'hC0; 15'h3AFA: d <= 8'hC0; 15'h3AFB: d <= 8'hC0;
                15'h3AFC: d <= 8'hC0; 15'h3AFD: d <= 8'hC0; 15'h3AFE: d <= 8'hC0; 15'h3AFF: d <= 8'hC0;
                15'h3B00: d <= 8'hC0; 15'h3B01: d <= 8'hC0; 15'h3B02: d <= 8'hC0; 15'h3B03: d <= 8'hC0;
                15'h3B04: d <= 8'hC0; 15'h3B05: d <= 8'hC0; 15'h3B06: d <= 8'hC0; 15'h3B07: d <= 8'hC0;
                15'h3B08: d <= 8'hC0; 15'h3B09: d <= 8'hC0; 15'h3B0A: d <= 8'hC0; 15'h3B0B: d <= 8'hC0;
                15'h3B0C: d <= 8'hC0; 15'h3B0D: d <= 8'hC0; 15'h3B0E: d <= 8'hC0; 15'h3B0F: d <= 8'hC0;
                15'h3B10: d <= 8'hC0; 15'h3B11: d <= 8'hC0; 15'h3B12: d <= 8'hC0; 15'h3B13: d <= 8'hC0;
                15'h3B14: d <= 8'hC0; 15'h3B15: d <= 8'hC0; 15'h3B16: d <= 8'hC0; 15'h3B17: d <= 8'hC0;
                15'h3B18: d <= 8'hC0; 15'h3B19: d <= 8'hC0; 15'h3B1A: d <= 8'hC0; 15'h3B1B: d <= 8'hC0;
                15'h3B1C: d <= 8'hC0; 15'h3B1D: d <= 8'hC0; 15'h3B1E: d <= 8'hC0; 15'h3B1F: d <= 8'hC0;
                15'h3B20: d <= 8'hC0; 15'h3B21: d <= 8'hC0; 15'h3B22: d <= 8'hC0; 15'h3B23: d <= 8'hC0;
                15'h3B24: d <= 8'hC0; 15'h3B25: d <= 8'hC0; 15'h3B26: d <= 8'hC0; 15'h3B27: d <= 8'hC0;
                15'h3B28: d <= 8'hC0; 15'h3B29: d <= 8'hC0; 15'h3B2A: d <= 8'hC0; 15'h3B2B: d <= 8'hC0;
                15'h3B2C: d <= 8'hC0; 15'h3B2D: d <= 8'hC0; 15'h3B2E: d <= 8'hC0; 15'h3B2F: d <= 8'hC0;
                15'h3B30: d <= 8'hC0; 15'h3B31: d <= 8'hC0; 15'h3B32: d <= 8'hC0; 15'h3B33: d <= 8'hC0;
                15'h3B34: d <= 8'hC0; 15'h3B35: d <= 8'hC0; 15'h3B36: d <= 8'hC0; 15'h3B37: d <= 8'hC0;
                15'h3B38: d <= 8'hC0; 15'h3B39: d <= 8'hC0; 15'h3B3A: d <= 8'hC0; 15'h3B3B: d <= 8'hC0;
                15'h3B3C: d <= 8'hC0; 15'h3B3D: d <= 8'hC0; 15'h3B3E: d <= 8'hC0; 15'h3B3F: d <= 8'hC0;
                15'h3B40: d <= 8'hC0; 15'h3B41: d <= 8'hC0; 15'h3B42: d <= 8'hC0; 15'h3B43: d <= 8'hC0;
                15'h3B44: d <= 8'hC0; 15'h3B45: d <= 8'hC0; 15'h3B46: d <= 8'hC0; 15'h3B47: d <= 8'hC0;
                15'h3B48: d <= 8'hC0; 15'h3B49: d <= 8'hC0; 15'h3B4A: d <= 8'hC0; 15'h3B4B: d <= 8'hC0;
                15'h3B4C: d <= 8'hC0; 15'h3B4D: d <= 8'hC0; 15'h3B4E: d <= 8'hC0; 15'h3B4F: d <= 8'hC0;
                15'h3B50: d <= 8'hC0; 15'h3B51: d <= 8'hC0; 15'h3B52: d <= 8'hC0; 15'h3B53: d <= 8'hC0;
                15'h3B54: d <= 8'hC0; 15'h3B55: d <= 8'hC0; 15'h3B56: d <= 8'hC0; 15'h3B57: d <= 8'hC0;
                15'h3B58: d <= 8'hC0; 15'h3B59: d <= 8'hC0; 15'h3B5A: d <= 8'hC0; 15'h3B5B: d <= 8'hC0;
                15'h3B5C: d <= 8'hC0; 15'h3B5D: d <= 8'hC0; 15'h3B5E: d <= 8'hC0; 15'h3B5F: d <= 8'hC0;
                15'h3B60: d <= 8'hC0; 15'h3B61: d <= 8'hC0; 15'h3B62: d <= 8'hC0; 15'h3B63: d <= 8'hC0;
                15'h3B64: d <= 8'hC0; 15'h3B65: d <= 8'hC0; 15'h3B66: d <= 8'hC0; 15'h3B67: d <= 8'hC0;
                15'h3B68: d <= 8'hC0; 15'h3B69: d <= 8'hC0; 15'h3B6A: d <= 8'hC0; 15'h3B6B: d <= 8'hC0;
                15'h3B6C: d <= 8'hC0; 15'h3B6D: d <= 8'hC0; 15'h3B6E: d <= 8'hC0; 15'h3B6F: d <= 8'hC0;
                15'h3B70: d <= 8'hC0; 15'h3B71: d <= 8'hC0; 15'h3B72: d <= 8'hC0; 15'h3B73: d <= 8'hC0;
                15'h3B74: d <= 8'hC0; 15'h3B75: d <= 8'hC0; 15'h3B76: d <= 8'hC0; 15'h3B77: d <= 8'hC0;
                15'h3B78: d <= 8'hC0; 15'h3B79: d <= 8'hC0; 15'h3B7A: d <= 8'hC0; 15'h3B7B: d <= 8'hC0;
                15'h3B7C: d <= 8'hC0; 15'h3B7D: d <= 8'hC0; 15'h3B7E: d <= 8'hC0; 15'h3B7F: d <= 8'hC0;
                15'h3B80: d <= 8'hC0; 15'h3B81: d <= 8'hC0; 15'h3B82: d <= 8'hC0; 15'h3B83: d <= 8'hC0;
                15'h3B84: d <= 8'hC0; 15'h3B85: d <= 8'hC0; 15'h3B86: d <= 8'hC0; 15'h3B87: d <= 8'hC0;
                15'h3B88: d <= 8'hC0; 15'h3B89: d <= 8'hC0; 15'h3B8A: d <= 8'hC0; 15'h3B8B: d <= 8'hC0;
                15'h3B8C: d <= 8'hC0; 15'h3B8D: d <= 8'hC0; 15'h3B8E: d <= 8'hC0; 15'h3B8F: d <= 8'hC0;
                15'h3B90: d <= 8'hC0; 15'h3B91: d <= 8'hC0; 15'h3B92: d <= 8'hC0; 15'h3B93: d <= 8'hC0;
                15'h3B94: d <= 8'hC0; 15'h3B95: d <= 8'hC0; 15'h3B96: d <= 8'hC0; 15'h3B97: d <= 8'hC0;
                15'h3B98: d <= 8'hC0; 15'h3B99: d <= 8'hC0; 15'h3B9A: d <= 8'hC0; 15'h3B9B: d <= 8'hC0;
                15'h3B9C: d <= 8'hC0; 15'h3B9D: d <= 8'hC0; 15'h3B9E: d <= 8'hC0; 15'h3B9F: d <= 8'hC0;
                15'h3BA0: d <= 8'hC0; 15'h3BA1: d <= 8'hC0; 15'h3BA2: d <= 8'hC0; 15'h3BA3: d <= 8'hC0;
                15'h3BA4: d <= 8'hC0; 15'h3BA5: d <= 8'hC0; 15'h3BA6: d <= 8'hC0; 15'h3BA7: d <= 8'hC0;
                15'h3BA8: d <= 8'hC0; 15'h3BA9: d <= 8'hC0; 15'h3BAA: d <= 8'hC0; 15'h3BAB: d <= 8'hC0;
                15'h3BAC: d <= 8'hC0; 15'h3BAD: d <= 8'hC0; 15'h3BAE: d <= 8'hC0; 15'h3BAF: d <= 8'hC0;
                15'h3BB0: d <= 8'hC0; 15'h3BB1: d <= 8'hC0; 15'h3BB2: d <= 8'hC0; 15'h3BB3: d <= 8'hC0;
                15'h3BB4: d <= 8'hC0; 15'h3BB5: d <= 8'hC0; 15'h3BB6: d <= 8'hC0; 15'h3BB7: d <= 8'hC0;
                15'h3BB8: d <= 8'hC0; 15'h3BB9: d <= 8'hC0; 15'h3BBA: d <= 8'hC0; 15'h3BBB: d <= 8'hC0;
                15'h3BBC: d <= 8'hC0; 15'h3BBD: d <= 8'hC0; 15'h3BBE: d <= 8'hC0; 15'h3BBF: d <= 8'hC0;
                15'h3BC0: d <= 8'hC0; 15'h3BC1: d <= 8'hC0; 15'h3BC2: d <= 8'hC0; 15'h3BC3: d <= 8'hC0;
                15'h3BC4: d <= 8'hC0; 15'h3BC5: d <= 8'hC0; 15'h3BC6: d <= 8'hC0; 15'h3BC7: d <= 8'hC0;
                15'h3BC8: d <= 8'hC0; 15'h3BC9: d <= 8'hC0; 15'h3BCA: d <= 8'hC0; 15'h3BCB: d <= 8'hC0;
                15'h3BCC: d <= 8'hC0; 15'h3BCD: d <= 8'hC0; 15'h3BCE: d <= 8'hC0; 15'h3BCF: d <= 8'hC0;
                15'h3BD0: d <= 8'hC0; 15'h3BD1: d <= 8'hC0; 15'h3BD2: d <= 8'hC0; 15'h3BD3: d <= 8'hC0;
                15'h3BD4: d <= 8'hC0; 15'h3BD5: d <= 8'hC0; 15'h3BD6: d <= 8'hC0; 15'h3BD7: d <= 8'hC0;
                15'h3BD8: d <= 8'hC0; 15'h3BD9: d <= 8'hC0; 15'h3BDA: d <= 8'hC0; 15'h3BDB: d <= 8'hC0;
                15'h3BDC: d <= 8'hC0; 15'h3BDD: d <= 8'hC0; 15'h3BDE: d <= 8'hC0; 15'h3BDF: d <= 8'hC0;
                15'h3BE0: d <= 8'hC0; 15'h3BE1: d <= 8'hC0; 15'h3BE2: d <= 8'hC0; 15'h3BE3: d <= 8'hC0;
                15'h3BE4: d <= 8'hC0; 15'h3BE5: d <= 8'hC0; 15'h3BE6: d <= 8'hC0; 15'h3BE7: d <= 8'hC0;
                15'h3BE8: d <= 8'hC0; 15'h3BE9: d <= 8'hC0; 15'h3BEA: d <= 8'hC0; 15'h3BEB: d <= 8'hC0;
                15'h3BEC: d <= 8'hC0; 15'h3BED: d <= 8'hC0; 15'h3BEE: d <= 8'hC0; 15'h3BEF: d <= 8'hC0;
                15'h3BF0: d <= 8'hC0; 15'h3BF1: d <= 8'hC0; 15'h3BF2: d <= 8'hC0; 15'h3BF3: d <= 8'hC0;
                15'h3BF4: d <= 8'hC0; 15'h3BF5: d <= 8'hC0; 15'h3BF6: d <= 8'hC0; 15'h3BF7: d <= 8'hC0;
                15'h3BF8: d <= 8'hC0; 15'h3BF9: d <= 8'hC0; 15'h3BFA: d <= 8'hC0; 15'h3BFB: d <= 8'hC0;
                15'h3BFC: d <= 8'hC0; 15'h3BFD: d <= 8'hC0; 15'h3BFE: d <= 8'hC0; 15'h3BFF: d <= 8'hC0;
                15'h3C00: d <= 8'hC0; 15'h3C01: d <= 8'hC0; 15'h3C02: d <= 8'hC0; 15'h3C03: d <= 8'hC0;
                15'h3C04: d <= 8'hC0; 15'h3C05: d <= 8'hC0; 15'h3C06: d <= 8'hC0; 15'h3C07: d <= 8'hC0;
                15'h3C08: d <= 8'hC0; 15'h3C09: d <= 8'hC0; 15'h3C0A: d <= 8'hC0; 15'h3C0B: d <= 8'hC0;
                15'h3C0C: d <= 8'hC0; 15'h3C0D: d <= 8'hC0; 15'h3C0E: d <= 8'hC0; 15'h3C0F: d <= 8'hC0;
                15'h3C10: d <= 8'hC0; 15'h3C11: d <= 8'hC0; 15'h3C12: d <= 8'hC0; 15'h3C13: d <= 8'hC0;
                15'h3C14: d <= 8'hC0; 15'h3C15: d <= 8'hC0; 15'h3C16: d <= 8'hC0; 15'h3C17: d <= 8'hC0;
                15'h3C18: d <= 8'hC0; 15'h3C19: d <= 8'hC0; 15'h3C1A: d <= 8'hC0; 15'h3C1B: d <= 8'hC0;
                15'h3C1C: d <= 8'hC0; 15'h3C1D: d <= 8'hC0; 15'h3C1E: d <= 8'hC0; 15'h3C1F: d <= 8'hC0;
                15'h3C20: d <= 8'hC0; 15'h3C21: d <= 8'hC0; 15'h3C22: d <= 8'hC0; 15'h3C23: d <= 8'hC0;
                15'h3C24: d <= 8'hC0; 15'h3C25: d <= 8'hC0; 15'h3C26: d <= 8'hC0; 15'h3C27: d <= 8'hC0;
                15'h3C28: d <= 8'hC0; 15'h3C29: d <= 8'hC0; 15'h3C2A: d <= 8'hC0; 15'h3C2B: d <= 8'hC0;
                15'h3C2C: d <= 8'hC0; 15'h3C2D: d <= 8'hC0; 15'h3C2E: d <= 8'hC0; 15'h3C2F: d <= 8'hC0;
                15'h3C30: d <= 8'hC0; 15'h3C31: d <= 8'hC0; 15'h3C32: d <= 8'hC0; 15'h3C33: d <= 8'hC0;
                15'h3C34: d <= 8'hC0; 15'h3C35: d <= 8'hC0; 15'h3C36: d <= 8'hC0; 15'h3C37: d <= 8'hC0;
                15'h3C38: d <= 8'hC0; 15'h3C39: d <= 8'hC0; 15'h3C3A: d <= 8'hC0; 15'h3C3B: d <= 8'hC0;
                15'h3C3C: d <= 8'hC0; 15'h3C3D: d <= 8'hC0; 15'h3C3E: d <= 8'hC0; 15'h3C3F: d <= 8'hC0;
                15'h3C40: d <= 8'hC0; 15'h3C41: d <= 8'hC0; 15'h3C42: d <= 8'hC0; 15'h3C43: d <= 8'hC0;
                15'h3C44: d <= 8'hC0; 15'h3C45: d <= 8'hC0; 15'h3C46: d <= 8'hC0; 15'h3C47: d <= 8'hC0;
                15'h3C48: d <= 8'hC0; 15'h3C49: d <= 8'hC0; 15'h3C4A: d <= 8'hC0; 15'h3C4B: d <= 8'hC0;
                15'h3C4C: d <= 8'hC0; 15'h3C4D: d <= 8'hC0; 15'h3C4E: d <= 8'hC0; 15'h3C4F: d <= 8'hC0;
                15'h3C50: d <= 8'hC0; 15'h3C51: d <= 8'hC0; 15'h3C52: d <= 8'hC0; 15'h3C53: d <= 8'hC0;
                15'h3C54: d <= 8'hC0; 15'h3C55: d <= 8'hC0; 15'h3C56: d <= 8'hC0; 15'h3C57: d <= 8'hC0;
                15'h3C58: d <= 8'hC0; 15'h3C59: d <= 8'hC0; 15'h3C5A: d <= 8'hC0; 15'h3C5B: d <= 8'hC0;
                15'h3C5C: d <= 8'hC0; 15'h3C5D: d <= 8'hC0; 15'h3C5E: d <= 8'hC0; 15'h3C5F: d <= 8'hC0;
                15'h3C60: d <= 8'hC0; 15'h3C61: d <= 8'hC0; 15'h3C62: d <= 8'hC0; 15'h3C63: d <= 8'hC0;
                15'h3C64: d <= 8'hC0; 15'h3C65: d <= 8'hC0; 15'h3C66: d <= 8'hC0; 15'h3C67: d <= 8'hC0;
                15'h3C68: d <= 8'hC0; 15'h3C69: d <= 8'hC0; 15'h3C6A: d <= 8'hC0; 15'h3C6B: d <= 8'hC0;
                15'h3C6C: d <= 8'hC0; 15'h3C6D: d <= 8'hC0; 15'h3C6E: d <= 8'hC0; 15'h3C6F: d <= 8'hC0;
                15'h3C70: d <= 8'hC0; 15'h3C71: d <= 8'hC0; 15'h3C72: d <= 8'hC0; 15'h3C73: d <= 8'hC0;
                15'h3C74: d <= 8'hC0; 15'h3C75: d <= 8'hC0; 15'h3C76: d <= 8'hC0; 15'h3C77: d <= 8'hC0;
                15'h3C78: d <= 8'hC0; 15'h3C79: d <= 8'hC0; 15'h3C7A: d <= 8'hC0; 15'h3C7B: d <= 8'hC0;
                15'h3C7C: d <= 8'hC0; 15'h3C7D: d <= 8'hC0; 15'h3C7E: d <= 8'hC0; 15'h3C7F: d <= 8'hC0;
                15'h3C80: d <= 8'hC0; 15'h3C81: d <= 8'hC0; 15'h3C82: d <= 8'hC0; 15'h3C83: d <= 8'hC0;
                15'h3C84: d <= 8'hC0; 15'h3C85: d <= 8'hC0; 15'h3C86: d <= 8'hC0; 15'h3C87: d <= 8'hC0;
                15'h3C88: d <= 8'hC0; 15'h3C89: d <= 8'hC0; 15'h3C8A: d <= 8'hC0; 15'h3C8B: d <= 8'hC0;
                15'h3C8C: d <= 8'hC0; 15'h3C8D: d <= 8'hC0; 15'h3C8E: d <= 8'hC0; 15'h3C8F: d <= 8'hC0;
                15'h3C90: d <= 8'hC0; 15'h3C91: d <= 8'hC0; 15'h3C92: d <= 8'hC0; 15'h3C93: d <= 8'hC0;
                15'h3C94: d <= 8'hC0; 15'h3C95: d <= 8'hC0; 15'h3C96: d <= 8'hC0; 15'h3C97: d <= 8'hC0;
                15'h3C98: d <= 8'hC0; 15'h3C99: d <= 8'hC0; 15'h3C9A: d <= 8'hC0; 15'h3C9B: d <= 8'hC0;
                15'h3C9C: d <= 8'hC0; 15'h3C9D: d <= 8'hC0; 15'h3C9E: d <= 8'hC0; 15'h3C9F: d <= 8'hC0;
                15'h3CA0: d <= 8'hC0; 15'h3CA1: d <= 8'hC0; 15'h3CA2: d <= 8'hC0; 15'h3CA3: d <= 8'hC0;
                15'h3CA4: d <= 8'hC0; 15'h3CA5: d <= 8'hC0; 15'h3CA6: d <= 8'hC0; 15'h3CA7: d <= 8'hC0;
                15'h3CA8: d <= 8'hC0; 15'h3CA9: d <= 8'hC0; 15'h3CAA: d <= 8'hC0; 15'h3CAB: d <= 8'hC0;
                15'h3CAC: d <= 8'hC0; 15'h3CAD: d <= 8'hC0; 15'h3CAE: d <= 8'hC0; 15'h3CAF: d <= 8'hC0;
                15'h3CB0: d <= 8'hC0; 15'h3CB1: d <= 8'hC0; 15'h3CB2: d <= 8'hC0; 15'h3CB3: d <= 8'hC0;
                15'h3CB4: d <= 8'hC0; 15'h3CB5: d <= 8'hC0; 15'h3CB6: d <= 8'hC0; 15'h3CB7: d <= 8'hC0;
                15'h3CB8: d <= 8'hC0; 15'h3CB9: d <= 8'hC0; 15'h3CBA: d <= 8'hC0; 15'h3CBB: d <= 8'hC0;
                15'h3CBC: d <= 8'hC0; 15'h3CBD: d <= 8'hC0; 15'h3CBE: d <= 8'hC0; 15'h3CBF: d <= 8'hC0;
                15'h3CC0: d <= 8'hC0; 15'h3CC1: d <= 8'hC0; 15'h3CC2: d <= 8'hC0; 15'h3CC3: d <= 8'hC0;
                15'h3CC4: d <= 8'hC0; 15'h3CC5: d <= 8'hC0; 15'h3CC6: d <= 8'hC0; 15'h3CC7: d <= 8'hC0;
                15'h3CC8: d <= 8'hC0; 15'h3CC9: d <= 8'hC0; 15'h3CCA: d <= 8'hC0; 15'h3CCB: d <= 8'hC0;
                15'h3CCC: d <= 8'hC0; 15'h3CCD: d <= 8'hC0; 15'h3CCE: d <= 8'hC0; 15'h3CCF: d <= 8'hC0;
                15'h3CD0: d <= 8'hC0; 15'h3CD1: d <= 8'hC0; 15'h3CD2: d <= 8'hC0; 15'h3CD3: d <= 8'hC0;
                15'h3CD4: d <= 8'hC0; 15'h3CD5: d <= 8'hC0; 15'h3CD6: d <= 8'hC0; 15'h3CD7: d <= 8'hC0;
                15'h3CD8: d <= 8'hC0; 15'h3CD9: d <= 8'hC0; 15'h3CDA: d <= 8'hC0; 15'h3CDB: d <= 8'hC0;
                15'h3CDC: d <= 8'hC0; 15'h3CDD: d <= 8'hC0; 15'h3CDE: d <= 8'hC0; 15'h3CDF: d <= 8'hC0;
                15'h3CE0: d <= 8'hC0; 15'h3CE1: d <= 8'hC0; 15'h3CE2: d <= 8'hC0; 15'h3CE3: d <= 8'hC0;
                15'h3CE4: d <= 8'hC0; 15'h3CE5: d <= 8'hC0; 15'h3CE6: d <= 8'hC0; 15'h3CE7: d <= 8'hC0;
                15'h3CE8: d <= 8'hC0; 15'h3CE9: d <= 8'hC0; 15'h3CEA: d <= 8'hC0; 15'h3CEB: d <= 8'hC0;
                15'h3CEC: d <= 8'hC0; 15'h3CED: d <= 8'hC0; 15'h3CEE: d <= 8'hC0; 15'h3CEF: d <= 8'hC0;
                15'h3CF0: d <= 8'hC0; 15'h3CF1: d <= 8'hC0; 15'h3CF2: d <= 8'hC0; 15'h3CF3: d <= 8'hC0;
                15'h3CF4: d <= 8'hC0; 15'h3CF5: d <= 8'hC0; 15'h3CF6: d <= 8'hC0; 15'h3CF7: d <= 8'hC0;
                15'h3CF8: d <= 8'hC0; 15'h3CF9: d <= 8'hC0; 15'h3CFA: d <= 8'hC0; 15'h3CFB: d <= 8'hC0;
                15'h3CFC: d <= 8'hC0; 15'h3CFD: d <= 8'hC0; 15'h3CFE: d <= 8'hC0; 15'h3CFF: d <= 8'hC0;
                15'h3D00: d <= 8'hC0; 15'h3D01: d <= 8'hC0; 15'h3D02: d <= 8'hC0; 15'h3D03: d <= 8'hC0;
                15'h3D04: d <= 8'hC0; 15'h3D05: d <= 8'hC0; 15'h3D06: d <= 8'hC0; 15'h3D07: d <= 8'hC0;
                15'h3D08: d <= 8'hC0; 15'h3D09: d <= 8'hC0; 15'h3D0A: d <= 8'hC0; 15'h3D0B: d <= 8'hC0;
                15'h3D0C: d <= 8'hC0; 15'h3D0D: d <= 8'hC0; 15'h3D0E: d <= 8'hC0; 15'h3D0F: d <= 8'hC0;
                15'h3D10: d <= 8'hC0; 15'h3D11: d <= 8'hC0; 15'h3D12: d <= 8'hC0; 15'h3D13: d <= 8'hC0;
                15'h3D14: d <= 8'hC0; 15'h3D15: d <= 8'hC0; 15'h3D16: d <= 8'hC0; 15'h3D17: d <= 8'hC0;
                15'h3D18: d <= 8'hC0; 15'h3D19: d <= 8'hC0; 15'h3D1A: d <= 8'hC0; 15'h3D1B: d <= 8'hC0;
                15'h3D1C: d <= 8'hC0; 15'h3D1D: d <= 8'hC0; 15'h3D1E: d <= 8'hC0; 15'h3D1F: d <= 8'hC0;
                15'h3D20: d <= 8'hC0; 15'h3D21: d <= 8'hC0; 15'h3D22: d <= 8'hC0; 15'h3D23: d <= 8'hC0;
                15'h3D24: d <= 8'hC0; 15'h3D25: d <= 8'hC0; 15'h3D26: d <= 8'hC0; 15'h3D27: d <= 8'hC0;
                15'h3D28: d <= 8'hC0; 15'h3D29: d <= 8'hC0; 15'h3D2A: d <= 8'hC0; 15'h3D2B: d <= 8'hC0;
                15'h3D2C: d <= 8'hC0; 15'h3D2D: d <= 8'hC0; 15'h3D2E: d <= 8'hC0; 15'h3D2F: d <= 8'hC0;
                15'h3D30: d <= 8'hC0; 15'h3D31: d <= 8'hC0; 15'h3D32: d <= 8'hC0; 15'h3D33: d <= 8'hC0;
                15'h3D34: d <= 8'hC0; 15'h3D35: d <= 8'hC0; 15'h3D36: d <= 8'hC0; 15'h3D37: d <= 8'hC0;
                15'h3D38: d <= 8'hC0; 15'h3D39: d <= 8'hC0; 15'h3D3A: d <= 8'hC0; 15'h3D3B: d <= 8'hC0;
                15'h3D3C: d <= 8'hC0; 15'h3D3D: d <= 8'hC0; 15'h3D3E: d <= 8'hC0; 15'h3D3F: d <= 8'hC0;
                15'h3D40: d <= 8'hC0; 15'h3D41: d <= 8'hC0; 15'h3D42: d <= 8'hC0; 15'h3D43: d <= 8'hC0;
                15'h3D44: d <= 8'hC0; 15'h3D45: d <= 8'hC0; 15'h3D46: d <= 8'hC0; 15'h3D47: d <= 8'hC0;
                15'h3D48: d <= 8'hC0; 15'h3D49: d <= 8'hC0; 15'h3D4A: d <= 8'hC0; 15'h3D4B: d <= 8'hC0;
                15'h3D4C: d <= 8'hC0; 15'h3D4D: d <= 8'hC0; 15'h3D4E: d <= 8'hC0; 15'h3D4F: d <= 8'hC0;
                15'h3D50: d <= 8'hC0; 15'h3D51: d <= 8'hC0; 15'h3D52: d <= 8'hC0; 15'h3D53: d <= 8'hC0;
                15'h3D54: d <= 8'hC0; 15'h3D55: d <= 8'hC0; 15'h3D56: d <= 8'hC0; 15'h3D57: d <= 8'hC0;
                15'h3D58: d <= 8'hC0; 15'h3D59: d <= 8'hC0; 15'h3D5A: d <= 8'hC0; 15'h3D5B: d <= 8'hC0;
                15'h3D5C: d <= 8'hC0; 15'h3D5D: d <= 8'hC0; 15'h3D5E: d <= 8'hC0; 15'h3D5F: d <= 8'hC0;
                15'h3D60: d <= 8'hC0; 15'h3D61: d <= 8'hC0; 15'h3D62: d <= 8'hC0; 15'h3D63: d <= 8'hC0;
                15'h3D64: d <= 8'hC0; 15'h3D65: d <= 8'hC0; 15'h3D66: d <= 8'hC0; 15'h3D67: d <= 8'hC0;
                15'h3D68: d <= 8'hC0; 15'h3D69: d <= 8'hC0; 15'h3D6A: d <= 8'hC0; 15'h3D6B: d <= 8'hC0;
                15'h3D6C: d <= 8'hC0; 15'h3D6D: d <= 8'hC0; 15'h3D6E: d <= 8'hC0; 15'h3D6F: d <= 8'hC0;
                15'h3D70: d <= 8'hC0; 15'h3D71: d <= 8'hC0; 15'h3D72: d <= 8'hC0; 15'h3D73: d <= 8'hC0;
                15'h3D74: d <= 8'hC0; 15'h3D75: d <= 8'hC0; 15'h3D76: d <= 8'hC0; 15'h3D77: d <= 8'hC0;
                15'h3D78: d <= 8'hC0; 15'h3D79: d <= 8'hC0; 15'h3D7A: d <= 8'hC0; 15'h3D7B: d <= 8'hC0;
                15'h3D7C: d <= 8'hC0; 15'h3D7D: d <= 8'hC0; 15'h3D7E: d <= 8'hC0; 15'h3D7F: d <= 8'hC0;
                15'h3D80: d <= 8'hC0; 15'h3D81: d <= 8'hC0; 15'h3D82: d <= 8'hC0; 15'h3D83: d <= 8'hC0;
                15'h3D84: d <= 8'hC0; 15'h3D85: d <= 8'hC0; 15'h3D86: d <= 8'hC0; 15'h3D87: d <= 8'hC0;
                15'h3D88: d <= 8'hC0; 15'h3D89: d <= 8'hC0; 15'h3D8A: d <= 8'hC0; 15'h3D8B: d <= 8'hC0;
                15'h3D8C: d <= 8'hC0; 15'h3D8D: d <= 8'hC0; 15'h3D8E: d <= 8'hC0; 15'h3D8F: d <= 8'hC0;
                15'h3D90: d <= 8'hC0; 15'h3D91: d <= 8'hC0; 15'h3D92: d <= 8'hC0; 15'h3D93: d <= 8'hC0;
                15'h3D94: d <= 8'hC0; 15'h3D95: d <= 8'hC0; 15'h3D96: d <= 8'hC0; 15'h3D97: d <= 8'hC0;
                15'h3D98: d <= 8'hC0; 15'h3D99: d <= 8'hC0; 15'h3D9A: d <= 8'hC0; 15'h3D9B: d <= 8'hC0;
                15'h3D9C: d <= 8'hC0; 15'h3D9D: d <= 8'hC0; 15'h3D9E: d <= 8'hC0; 15'h3D9F: d <= 8'hC0;
                15'h3DA0: d <= 8'hC0; 15'h3DA1: d <= 8'hC0; 15'h3DA2: d <= 8'hC0; 15'h3DA3: d <= 8'hC0;
                15'h3DA4: d <= 8'hC0; 15'h3DA5: d <= 8'hC0; 15'h3DA6: d <= 8'hC0; 15'h3DA7: d <= 8'hC0;
                15'h3DA8: d <= 8'hC0; 15'h3DA9: d <= 8'hC0; 15'h3DAA: d <= 8'hC0; 15'h3DAB: d <= 8'hC0;
                15'h3DAC: d <= 8'hC0; 15'h3DAD: d <= 8'hC0; 15'h3DAE: d <= 8'hC0; 15'h3DAF: d <= 8'hC0;
                15'h3DB0: d <= 8'hC0; 15'h3DB1: d <= 8'hC0; 15'h3DB2: d <= 8'hC0; 15'h3DB3: d <= 8'hC0;
                15'h3DB4: d <= 8'hC0; 15'h3DB5: d <= 8'hC0; 15'h3DB6: d <= 8'hC0; 15'h3DB7: d <= 8'hC0;
                15'h3DB8: d <= 8'hC0; 15'h3DB9: d <= 8'hC0; 15'h3DBA: d <= 8'hC0; 15'h3DBB: d <= 8'hC0;
                15'h3DBC: d <= 8'hC0; 15'h3DBD: d <= 8'hC0; 15'h3DBE: d <= 8'hC0; 15'h3DBF: d <= 8'hC0;
                15'h3DC0: d <= 8'hC0; 15'h3DC1: d <= 8'hC0; 15'h3DC2: d <= 8'hC0; 15'h3DC3: d <= 8'hC0;
                15'h3DC4: d <= 8'hC0; 15'h3DC5: d <= 8'hC0; 15'h3DC6: d <= 8'hC0; 15'h3DC7: d <= 8'hC0;
                15'h3DC8: d <= 8'hC0; 15'h3DC9: d <= 8'hC0; 15'h3DCA: d <= 8'hC0; 15'h3DCB: d <= 8'hC0;
                15'h3DCC: d <= 8'hC0; 15'h3DCD: d <= 8'hC0; 15'h3DCE: d <= 8'hC0; 15'h3DCF: d <= 8'hC0;
                15'h3DD0: d <= 8'hC0; 15'h3DD1: d <= 8'hC0; 15'h3DD2: d <= 8'hC0; 15'h3DD3: d <= 8'hC0;
                15'h3DD4: d <= 8'hC0; 15'h3DD5: d <= 8'hC0; 15'h3DD6: d <= 8'hC0; 15'h3DD7: d <= 8'hC0;
                15'h3DD8: d <= 8'hC0; 15'h3DD9: d <= 8'hC0; 15'h3DDA: d <= 8'hC0; 15'h3DDB: d <= 8'hC0;
                15'h3DDC: d <= 8'hC0; 15'h3DDD: d <= 8'hC0; 15'h3DDE: d <= 8'hC0; 15'h3DDF: d <= 8'hC0;
                15'h3DE0: d <= 8'hC0; 15'h3DE1: d <= 8'hC0; 15'h3DE2: d <= 8'hC0; 15'h3DE3: d <= 8'hC0;
                15'h3DE4: d <= 8'hC0; 15'h3DE5: d <= 8'hC0; 15'h3DE6: d <= 8'hC0; 15'h3DE7: d <= 8'hC0;
                15'h3DE8: d <= 8'hC0; 15'h3DE9: d <= 8'hC0; 15'h3DEA: d <= 8'hC0; 15'h3DEB: d <= 8'hC0;
                15'h3DEC: d <= 8'hC0; 15'h3DED: d <= 8'hC0; 15'h3DEE: d <= 8'hC0; 15'h3DEF: d <= 8'hC0;
                15'h3DF0: d <= 8'hC0; 15'h3DF1: d <= 8'hC0; 15'h3DF2: d <= 8'hC0; 15'h3DF3: d <= 8'hC0;
                15'h3DF4: d <= 8'hC0; 15'h3DF5: d <= 8'hC0; 15'h3DF6: d <= 8'hC0; 15'h3DF7: d <= 8'hC0;
                15'h3DF8: d <= 8'hC0; 15'h3DF9: d <= 8'hC0; 15'h3DFA: d <= 8'hC0; 15'h3DFB: d <= 8'hC0;
                15'h3DFC: d <= 8'hC0; 15'h3DFD: d <= 8'hC0; 15'h3DFE: d <= 8'hC0; 15'h3DFF: d <= 8'hC0;
                15'h3E00: d <= 8'hC0; 15'h3E01: d <= 8'hC0; 15'h3E02: d <= 8'hC0; 15'h3E03: d <= 8'hC0;
                15'h3E04: d <= 8'hC0; 15'h3E05: d <= 8'hC0; 15'h3E06: d <= 8'hC0; 15'h3E07: d <= 8'hC0;
                15'h3E08: d <= 8'hC0; 15'h3E09: d <= 8'hC0; 15'h3E0A: d <= 8'hC0; 15'h3E0B: d <= 8'hC0;
                15'h3E0C: d <= 8'hC0; 15'h3E0D: d <= 8'hC0; 15'h3E0E: d <= 8'hC0; 15'h3E0F: d <= 8'hC0;
                15'h3E10: d <= 8'hC0; 15'h3E11: d <= 8'hC0; 15'h3E12: d <= 8'hC0; 15'h3E13: d <= 8'hC0;
                15'h3E14: d <= 8'hC0; 15'h3E15: d <= 8'hC0; 15'h3E16: d <= 8'hC0; 15'h3E17: d <= 8'hC0;
                15'h3E18: d <= 8'hC0; 15'h3E19: d <= 8'hC0; 15'h3E1A: d <= 8'hC0; 15'h3E1B: d <= 8'hC0;
                15'h3E1C: d <= 8'hC0; 15'h3E1D: d <= 8'hC0; 15'h3E1E: d <= 8'hC0; 15'h3E1F: d <= 8'hC0;
                15'h3E20: d <= 8'hC0; 15'h3E21: d <= 8'hC0; 15'h3E22: d <= 8'hC0; 15'h3E23: d <= 8'hC0;
                15'h3E24: d <= 8'hC0; 15'h3E25: d <= 8'hC0; 15'h3E26: d <= 8'hC0; 15'h3E27: d <= 8'hC0;
                15'h3E28: d <= 8'hC0; 15'h3E29: d <= 8'hC0; 15'h3E2A: d <= 8'hC0; 15'h3E2B: d <= 8'hC0;
                15'h3E2C: d <= 8'hC0; 15'h3E2D: d <= 8'hC0; 15'h3E2E: d <= 8'hC0; 15'h3E2F: d <= 8'hC0;
                15'h3E30: d <= 8'hC0; 15'h3E31: d <= 8'hC0; 15'h3E32: d <= 8'hC0; 15'h3E33: d <= 8'hC0;
                15'h3E34: d <= 8'hC0; 15'h3E35: d <= 8'hC0; 15'h3E36: d <= 8'hC0; 15'h3E37: d <= 8'hC0;
                15'h3E38: d <= 8'hC0; 15'h3E39: d <= 8'hC0; 15'h3E3A: d <= 8'hC0; 15'h3E3B: d <= 8'hC0;
                15'h3E3C: d <= 8'hC0; 15'h3E3D: d <= 8'hC0; 15'h3E3E: d <= 8'hC0; 15'h3E3F: d <= 8'hC0;
                15'h3E40: d <= 8'hC0; 15'h3E41: d <= 8'hC0; 15'h3E42: d <= 8'hC0; 15'h3E43: d <= 8'hC0;
                15'h3E44: d <= 8'hC0; 15'h3E45: d <= 8'hC0; 15'h3E46: d <= 8'hC0; 15'h3E47: d <= 8'hC0;
                15'h3E48: d <= 8'hC0; 15'h3E49: d <= 8'hC0; 15'h3E4A: d <= 8'hC0; 15'h3E4B: d <= 8'hC0;
                15'h3E4C: d <= 8'hC0; 15'h3E4D: d <= 8'hC0; 15'h3E4E: d <= 8'hC0; 15'h3E4F: d <= 8'hC0;
                15'h3E50: d <= 8'hC0; 15'h3E51: d <= 8'hC0; 15'h3E52: d <= 8'hC0; 15'h3E53: d <= 8'hC0;
                15'h3E54: d <= 8'hC0; 15'h3E55: d <= 8'hC0; 15'h3E56: d <= 8'hC0; 15'h3E57: d <= 8'hC0;
                15'h3E58: d <= 8'hC0; 15'h3E59: d <= 8'hC0; 15'h3E5A: d <= 8'hC0; 15'h3E5B: d <= 8'hC0;
                15'h3E5C: d <= 8'hC0; 15'h3E5D: d <= 8'hC0; 15'h3E5E: d <= 8'hC0; 15'h3E5F: d <= 8'hC0;
                15'h3E60: d <= 8'hC0; 15'h3E61: d <= 8'hC0; 15'h3E62: d <= 8'hC0; 15'h3E63: d <= 8'hC0;
                15'h3E64: d <= 8'hC0; 15'h3E65: d <= 8'hC0; 15'h3E66: d <= 8'hC0; 15'h3E67: d <= 8'hC0;
                15'h3E68: d <= 8'hC0; 15'h3E69: d <= 8'hC0; 15'h3E6A: d <= 8'hC0; 15'h3E6B: d <= 8'hC0;
                15'h3E6C: d <= 8'hC0; 15'h3E6D: d <= 8'hC0; 15'h3E6E: d <= 8'hC0; 15'h3E6F: d <= 8'hC0;
                15'h3E70: d <= 8'hC0; 15'h3E71: d <= 8'hC0; 15'h3E72: d <= 8'hC0; 15'h3E73: d <= 8'hC0;
                15'h3E74: d <= 8'hC0; 15'h3E75: d <= 8'hC0; 15'h3E76: d <= 8'hC0; 15'h3E77: d <= 8'hC0;
                15'h3E78: d <= 8'hC0; 15'h3E79: d <= 8'hC0; 15'h3E7A: d <= 8'hC0; 15'h3E7B: d <= 8'hC0;
                15'h3E7C: d <= 8'hC0; 15'h3E7D: d <= 8'hC0; 15'h3E7E: d <= 8'hC0; 15'h3E7F: d <= 8'hC0;
                15'h3E80: d <= 8'hC0; 15'h3E81: d <= 8'hC0; 15'h3E82: d <= 8'hC0; 15'h3E83: d <= 8'hC0;
                15'h3E84: d <= 8'hC0; 15'h3E85: d <= 8'hC0; 15'h3E86: d <= 8'hC0; 15'h3E87: d <= 8'hC0;
                15'h3E88: d <= 8'hC0; 15'h3E89: d <= 8'hC0; 15'h3E8A: d <= 8'hC0; 15'h3E8B: d <= 8'hC0;
                15'h3E8C: d <= 8'hC0; 15'h3E8D: d <= 8'hC0; 15'h3E8E: d <= 8'hC0; 15'h3E8F: d <= 8'hC0;
                15'h3E90: d <= 8'hC0; 15'h3E91: d <= 8'hC0; 15'h3E92: d <= 8'hC0; 15'h3E93: d <= 8'hC0;
                15'h3E94: d <= 8'hC0; 15'h3E95: d <= 8'hC0; 15'h3E96: d <= 8'hC0; 15'h3E97: d <= 8'hC0;
                15'h3E98: d <= 8'hC0; 15'h3E99: d <= 8'hC0; 15'h3E9A: d <= 8'hC0; 15'h3E9B: d <= 8'hC0;
                15'h3E9C: d <= 8'hC0; 15'h3E9D: d <= 8'hC0; 15'h3E9E: d <= 8'hC0; 15'h3E9F: d <= 8'hC0;
                15'h3EA0: d <= 8'hC0; 15'h3EA1: d <= 8'hC0; 15'h3EA2: d <= 8'hC0; 15'h3EA3: d <= 8'hC0;
                15'h3EA4: d <= 8'hC0; 15'h3EA5: d <= 8'hC0; 15'h3EA6: d <= 8'hC0; 15'h3EA7: d <= 8'hC0;
                15'h3EA8: d <= 8'hC0; 15'h3EA9: d <= 8'hC0; 15'h3EAA: d <= 8'hC0; 15'h3EAB: d <= 8'hC0;
                15'h3EAC: d <= 8'hC0; 15'h3EAD: d <= 8'hC0; 15'h3EAE: d <= 8'hC0; 15'h3EAF: d <= 8'hC0;
                15'h3EB0: d <= 8'hC0; 15'h3EB1: d <= 8'hC0; 15'h3EB2: d <= 8'hC0; 15'h3EB3: d <= 8'hC0;
                15'h3EB4: d <= 8'hC0; 15'h3EB5: d <= 8'hC0; 15'h3EB6: d <= 8'hC0; 15'h3EB7: d <= 8'hC0;
                15'h3EB8: d <= 8'hC0; 15'h3EB9: d <= 8'hC0; 15'h3EBA: d <= 8'hC0; 15'h3EBB: d <= 8'hC0;
                15'h3EBC: d <= 8'hC0; 15'h3EBD: d <= 8'hC0; 15'h3EBE: d <= 8'hC0; 15'h3EBF: d <= 8'hC0;
                15'h3EC0: d <= 8'hC0; 15'h3EC1: d <= 8'hC0; 15'h3EC2: d <= 8'hC0; 15'h3EC3: d <= 8'hC0;
                15'h3EC4: d <= 8'hC0; 15'h3EC5: d <= 8'hC0; 15'h3EC6: d <= 8'hC0; 15'h3EC7: d <= 8'hC0;
                15'h3EC8: d <= 8'hC0; 15'h3EC9: d <= 8'hC0; 15'h3ECA: d <= 8'hC0; 15'h3ECB: d <= 8'hC0;
                15'h3ECC: d <= 8'hC0; 15'h3ECD: d <= 8'hC0; 15'h3ECE: d <= 8'hC0; 15'h3ECF: d <= 8'hC0;
                15'h3ED0: d <= 8'hC0; 15'h3ED1: d <= 8'hC0; 15'h3ED2: d <= 8'hC0; 15'h3ED3: d <= 8'hC0;
                15'h3ED4: d <= 8'hC0; 15'h3ED5: d <= 8'hC0; 15'h3ED6: d <= 8'hC0; 15'h3ED7: d <= 8'hC0;
                15'h3ED8: d <= 8'hC0; 15'h3ED9: d <= 8'hC0; 15'h3EDA: d <= 8'hC0; 15'h3EDB: d <= 8'hC0;
                15'h3EDC: d <= 8'hC0; 15'h3EDD: d <= 8'hC0; 15'h3EDE: d <= 8'hC0; 15'h3EDF: d <= 8'hC0;
                15'h3EE0: d <= 8'hC0; 15'h3EE1: d <= 8'hC0; 15'h3EE2: d <= 8'hC0; 15'h3EE3: d <= 8'hC0;
                15'h3EE4: d <= 8'hC0; 15'h3EE5: d <= 8'hC0; 15'h3EE6: d <= 8'hC0; 15'h3EE7: d <= 8'hC0;
                15'h3EE8: d <= 8'hC0; 15'h3EE9: d <= 8'hC0; 15'h3EEA: d <= 8'hC0; 15'h3EEB: d <= 8'hC0;
                15'h3EEC: d <= 8'hC0; 15'h3EED: d <= 8'hC0; 15'h3EEE: d <= 8'hC0; 15'h3EEF: d <= 8'hC0;
                15'h3EF0: d <= 8'hC0; 15'h3EF1: d <= 8'hC0; 15'h3EF2: d <= 8'hC0; 15'h3EF3: d <= 8'hC0;
                15'h3EF4: d <= 8'hC0; 15'h3EF5: d <= 8'hC0; 15'h3EF6: d <= 8'hC0; 15'h3EF7: d <= 8'hC0;
                15'h3EF8: d <= 8'hC0; 15'h3EF9: d <= 8'hC0; 15'h3EFA: d <= 8'hC0; 15'h3EFB: d <= 8'hC0;
                15'h3EFC: d <= 8'hC0; 15'h3EFD: d <= 8'hC0; 15'h3EFE: d <= 8'hC0; 15'h3EFF: d <= 8'hC0;
                15'h3F00: d <= 8'hC0; 15'h3F01: d <= 8'hC0; 15'h3F02: d <= 8'hC0; 15'h3F03: d <= 8'hC0;
                15'h3F04: d <= 8'hC0; 15'h3F05: d <= 8'hC0; 15'h3F06: d <= 8'hC0; 15'h3F07: d <= 8'hC0;
                15'h3F08: d <= 8'hC0; 15'h3F09: d <= 8'hC0; 15'h3F0A: d <= 8'hC0; 15'h3F0B: d <= 8'hC0;
                15'h3F0C: d <= 8'hC0; 15'h3F0D: d <= 8'hC0; 15'h3F0E: d <= 8'hC0; 15'h3F0F: d <= 8'hC0;
                15'h3F10: d <= 8'hC0; 15'h3F11: d <= 8'hC0; 15'h3F12: d <= 8'hC0; 15'h3F13: d <= 8'hC0;
                15'h3F14: d <= 8'hC0; 15'h3F15: d <= 8'hC0; 15'h3F16: d <= 8'hC0; 15'h3F17: d <= 8'hC0;
                15'h3F18: d <= 8'hC0; 15'h3F19: d <= 8'hC0; 15'h3F1A: d <= 8'hC0; 15'h3F1B: d <= 8'hC0;
                15'h3F1C: d <= 8'hC0; 15'h3F1D: d <= 8'hC0; 15'h3F1E: d <= 8'hC0; 15'h3F1F: d <= 8'hC0;
                15'h3F20: d <= 8'hC0; 15'h3F21: d <= 8'hC0; 15'h3F22: d <= 8'hC0; 15'h3F23: d <= 8'hC0;
                15'h3F24: d <= 8'hC0; 15'h3F25: d <= 8'hC0; 15'h3F26: d <= 8'hC0; 15'h3F27: d <= 8'hC0;
                15'h3F28: d <= 8'hC0; 15'h3F29: d <= 8'hC0; 15'h3F2A: d <= 8'hC0; 15'h3F2B: d <= 8'hC0;
                15'h3F2C: d <= 8'hC0; 15'h3F2D: d <= 8'hC0; 15'h3F2E: d <= 8'hC0; 15'h3F2F: d <= 8'hC0;
                15'h3F30: d <= 8'hC0; 15'h3F31: d <= 8'hC0; 15'h3F32: d <= 8'hC0; 15'h3F33: d <= 8'hC0;
                15'h3F34: d <= 8'hC0; 15'h3F35: d <= 8'hC0; 15'h3F36: d <= 8'hC0; 15'h3F37: d <= 8'hC0;
                15'h3F38: d <= 8'hC0; 15'h3F39: d <= 8'hC0; 15'h3F3A: d <= 8'hC0; 15'h3F3B: d <= 8'hC0;
                15'h3F3C: d <= 8'hC0; 15'h3F3D: d <= 8'hC0; 15'h3F3E: d <= 8'hC0; 15'h3F3F: d <= 8'hC0;
                15'h3F40: d <= 8'hC0; 15'h3F41: d <= 8'hC0; 15'h3F42: d <= 8'hC0; 15'h3F43: d <= 8'hC0;
                15'h3F44: d <= 8'hC0; 15'h3F45: d <= 8'hC0; 15'h3F46: d <= 8'hC0; 15'h3F47: d <= 8'hC0;
                15'h3F48: d <= 8'hC0; 15'h3F49: d <= 8'hC0; 15'h3F4A: d <= 8'hC0; 15'h3F4B: d <= 8'hC0;
                15'h3F4C: d <= 8'hC0; 15'h3F4D: d <= 8'hC0; 15'h3F4E: d <= 8'hC0; 15'h3F4F: d <= 8'hC0;
                15'h3F50: d <= 8'hC0; 15'h3F51: d <= 8'hC0; 15'h3F52: d <= 8'hC0; 15'h3F53: d <= 8'hC0;
                15'h3F54: d <= 8'hC0; 15'h3F55: d <= 8'hC0; 15'h3F56: d <= 8'hC0; 15'h3F57: d <= 8'hC0;
                15'h3F58: d <= 8'hC0; 15'h3F59: d <= 8'hC0; 15'h3F5A: d <= 8'hC0; 15'h3F5B: d <= 8'hC0;
                15'h3F5C: d <= 8'hC0; 15'h3F5D: d <= 8'hC0; 15'h3F5E: d <= 8'hC0; 15'h3F5F: d <= 8'hC0;
                15'h3F60: d <= 8'hC0; 15'h3F61: d <= 8'hC0; 15'h3F62: d <= 8'hC0; 15'h3F63: d <= 8'hC0;
                15'h3F64: d <= 8'hC0; 15'h3F65: d <= 8'hC0; 15'h3F66: d <= 8'hC0; 15'h3F67: d <= 8'hC0;
                15'h3F68: d <= 8'hC0; 15'h3F69: d <= 8'hC0; 15'h3F6A: d <= 8'hC0; 15'h3F6B: d <= 8'hC0;
                15'h3F6C: d <= 8'hC0; 15'h3F6D: d <= 8'hC0; 15'h3F6E: d <= 8'hC0; 15'h3F6F: d <= 8'hC0;
                15'h3F70: d <= 8'hC0; 15'h3F71: d <= 8'hC0; 15'h3F72: d <= 8'hC0; 15'h3F73: d <= 8'hC0;
                15'h3F74: d <= 8'hC0; 15'h3F75: d <= 8'hC0; 15'h3F76: d <= 8'hC0; 15'h3F77: d <= 8'hC0;
                15'h3F78: d <= 8'hC0; 15'h3F79: d <= 8'hC0; 15'h3F7A: d <= 8'hC0; 15'h3F7B: d <= 8'hC0;
                15'h3F7C: d <= 8'hC0; 15'h3F7D: d <= 8'hC0; 15'h3F7E: d <= 8'hC0; 15'h3F7F: d <= 8'hC0;
                15'h3F80: d <= 8'hC0; 15'h3F81: d <= 8'hC0; 15'h3F82: d <= 8'hC0; 15'h3F83: d <= 8'hC0;
                15'h3F84: d <= 8'hC0; 15'h3F85: d <= 8'hC0; 15'h3F86: d <= 8'hC0; 15'h3F87: d <= 8'hC0;
                15'h3F88: d <= 8'hC0; 15'h3F89: d <= 8'hC0; 15'h3F8A: d <= 8'hC0; 15'h3F8B: d <= 8'hC0;
                15'h3F8C: d <= 8'hC0; 15'h3F8D: d <= 8'hC0; 15'h3F8E: d <= 8'hC0; 15'h3F8F: d <= 8'hC0;
                15'h3F90: d <= 8'hC0; 15'h3F91: d <= 8'hC0; 15'h3F92: d <= 8'hC0; 15'h3F93: d <= 8'hC0;
                15'h3F94: d <= 8'hC0; 15'h3F95: d <= 8'hC0; 15'h3F96: d <= 8'hC0; 15'h3F97: d <= 8'hC0;
                15'h3F98: d <= 8'hC0; 15'h3F99: d <= 8'hC0; 15'h3F9A: d <= 8'hC0; 15'h3F9B: d <= 8'hC0;
                15'h3F9C: d <= 8'hC0; 15'h3F9D: d <= 8'hC0; 15'h3F9E: d <= 8'hC0; 15'h3F9F: d <= 8'hC0;
                15'h3FA0: d <= 8'hC0; 15'h3FA1: d <= 8'hC0; 15'h3FA2: d <= 8'hC0; 15'h3FA3: d <= 8'hC0;
                15'h3FA4: d <= 8'hC0; 15'h3FA5: d <= 8'hC0; 15'h3FA6: d <= 8'hC0; 15'h3FA7: d <= 8'hC0;
                15'h3FA8: d <= 8'hC0; 15'h3FA9: d <= 8'hC0; 15'h3FAA: d <= 8'hC0; 15'h3FAB: d <= 8'hC0;
                15'h3FAC: d <= 8'hC0; 15'h3FAD: d <= 8'hC0; 15'h3FAE: d <= 8'hC0; 15'h3FAF: d <= 8'hC0;
                15'h3FB0: d <= 8'hC0; 15'h3FB1: d <= 8'hC0; 15'h3FB2: d <= 8'hC0; 15'h3FB3: d <= 8'hC0;
                15'h3FB4: d <= 8'hC0; 15'h3FB5: d <= 8'hC0; 15'h3FB6: d <= 8'hC0; 15'h3FB7: d <= 8'hC0;
                15'h3FB8: d <= 8'hC0; 15'h3FB9: d <= 8'hC0; 15'h3FBA: d <= 8'hC0; 15'h3FBB: d <= 8'hC0;
                15'h3FBC: d <= 8'hC0; 15'h3FBD: d <= 8'hC0; 15'h3FBE: d <= 8'hC0; 15'h3FBF: d <= 8'hC0;
                15'h3FC0: d <= 8'hC0; 15'h3FC1: d <= 8'hC0; 15'h3FC2: d <= 8'hC0; 15'h3FC3: d <= 8'hC0;
                15'h3FC4: d <= 8'hC0; 15'h3FC5: d <= 8'hC0; 15'h3FC6: d <= 8'hC0; 15'h3FC7: d <= 8'hC0;
                15'h3FC8: d <= 8'hC0; 15'h3FC9: d <= 8'hC0; 15'h3FCA: d <= 8'hC0; 15'h3FCB: d <= 8'hC0;
                15'h3FCC: d <= 8'hC0; 15'h3FCD: d <= 8'hC0; 15'h3FCE: d <= 8'hC0; 15'h3FCF: d <= 8'hC0;
                15'h3FD0: d <= 8'hC0; 15'h3FD1: d <= 8'hC0; 15'h3FD2: d <= 8'hC0; 15'h3FD3: d <= 8'hC0;
                15'h3FD4: d <= 8'hC0; 15'h3FD5: d <= 8'hC0; 15'h3FD6: d <= 8'hC0; 15'h3FD7: d <= 8'hC0;
                15'h3FD8: d <= 8'hC0; 15'h3FD9: d <= 8'hC0; 15'h3FDA: d <= 8'hC0; 15'h3FDB: d <= 8'hC0;
                15'h3FDC: d <= 8'hC0; 15'h3FDD: d <= 8'hC0; 15'h3FDE: d <= 8'hC0; 15'h3FDF: d <= 8'hC0;
                15'h3FE0: d <= 8'hC0; 15'h3FE1: d <= 8'hC0; 15'h3FE2: d <= 8'hC0; 15'h3FE3: d <= 8'hC0;
                15'h3FE4: d <= 8'hC0; 15'h3FE5: d <= 8'hC0; 15'h3FE6: d <= 8'hC0; 15'h3FE7: d <= 8'hC0;
                15'h3FE8: d <= 8'hC0; 15'h3FE9: d <= 8'hC0; 15'h3FEA: d <= 8'hC0; 15'h3FEB: d <= 8'hC0;
                15'h3FEC: d <= 8'hC0; 15'h3FED: d <= 8'hC0; 15'h3FEE: d <= 8'hC0; 15'h3FEF: d <= 8'hC0;
                15'h3FF0: d <= 8'hC0; 15'h3FF1: d <= 8'hC0; 15'h3FF2: d <= 8'hC0; 15'h3FF3: d <= 8'hC0;
                15'h3FF4: d <= 8'hC0; 15'h3FF5: d <= 8'hC0; 15'h3FF6: d <= 8'hC0; 15'h3FF7: d <= 8'hC0;
                15'h3FF8: d <= 8'hC0; 15'h3FF9: d <= 8'hC0; 15'h3FFA: d <= 8'hC0; 15'h3FFB: d <= 8'hC0;
                15'h3FFC: d <= 8'hC0; 15'h3FFD: d <= 8'hC0; 15'h3FFE: d <= 8'hC0; 15'h3FFF: d <= 8'hC0;
                15'h4000: d <= 8'h00; 15'h4001: d <= 8'h00; 15'h4002: d <= 8'h00; 15'h4003: d <= 8'h00;
                15'h4004: d <= 8'h00; 15'h4005: d <= 8'h00; 15'h4006: d <= 8'h00; 15'h4007: d <= 8'h00;
                15'h4008: d <= 8'h00; 15'h4009: d <= 8'h00; 15'h400A: d <= 8'h00; 15'h400B: d <= 8'h00;
                15'h400C: d <= 8'h00; 15'h400D: d <= 8'h00; 15'h400E: d <= 8'h00; 15'h400F: d <= 8'h00;
                15'h4010: d <= 8'h00; 15'h4011: d <= 8'h00; 15'h4012: d <= 8'h00; 15'h4013: d <= 8'h00;
                15'h4014: d <= 8'h00; 15'h4015: d <= 8'h00; 15'h4016: d <= 8'h00; 15'h4017: d <= 8'h00;
                15'h4018: d <= 8'h00; 15'h4019: d <= 8'h00; 15'h401A: d <= 8'h00; 15'h401B: d <= 8'h00;
                15'h401C: d <= 8'h00; 15'h401D: d <= 8'h00; 15'h401E: d <= 8'h00; 15'h401F: d <= 8'h00;
                15'h4020: d <= 8'h00; 15'h4021: d <= 8'h00; 15'h4022: d <= 8'h00; 15'h4023: d <= 8'h00;
                15'h4024: d <= 8'h00; 15'h4025: d <= 8'h00; 15'h4026: d <= 8'h00; 15'h4027: d <= 8'h00;
                15'h4028: d <= 8'h00; 15'h4029: d <= 8'h00; 15'h402A: d <= 8'h00; 15'h402B: d <= 8'h00;
                15'h402C: d <= 8'h00; 15'h402D: d <= 8'h00; 15'h402E: d <= 8'h00; 15'h402F: d <= 8'hAF;
                15'h4030: d <= 8'h00; 15'h4031: d <= 8'h00; 15'h4032: d <= 8'h00; 15'h4033: d <= 8'h00;
                15'h4034: d <= 8'h00; 15'h4035: d <= 8'h00; 15'h4036: d <= 8'h00; 15'h4037: d <= 8'h00;
                15'h4038: d <= 8'h00; 15'h4039: d <= 8'h00; 15'h403A: d <= 8'h00; 15'h403B: d <= 8'h00;
                15'h403C: d <= 8'h00; 15'h403D: d <= 8'h00; 15'h403E: d <= 8'h00; 15'h403F: d <= 8'h00;
                15'h4040: d <= 8'h00; 15'h4041: d <= 8'h00; 15'h4042: d <= 8'h00; 15'h4043: d <= 8'h00;
                15'h4044: d <= 8'h00; 15'h4045: d <= 8'h00; 15'h4046: d <= 8'h00; 15'h4047: d <= 8'h00;
                15'h4048: d <= 8'h00; 15'h4049: d <= 8'h00; 15'h404A: d <= 8'h00; 15'h404B: d <= 8'h00;
                15'h404C: d <= 8'h00; 15'h404D: d <= 8'h00; 15'h404E: d <= 8'h00; 15'h404F: d <= 8'h00;
                15'h4050: d <= 8'h00; 15'h4051: d <= 8'h00; 15'h4052: d <= 8'h00; 15'h4053: d <= 8'h00;
                15'h4054: d <= 8'h00; 15'h4055: d <= 8'h00; 15'h4056: d <= 8'h00; 15'h4057: d <= 8'h00;
                15'h4058: d <= 8'h45; 15'h4059: d <= 8'h35; 15'h405A: d <= 8'hAA; 15'h405B: d <= 8'h00;
                15'h405C: d <= 8'h00; 15'h405D: d <= 8'h00; 15'h405E: d <= 8'h00; 15'h405F: d <= 8'h00;
                15'h4060: d <= 8'h00; 15'h4061: d <= 8'h00; 15'h4062: d <= 8'h00; 15'h4063: d <= 8'h00;
                15'h4064: d <= 8'h00; 15'h4065: d <= 8'h00; 15'h4066: d <= 8'h00; 15'h4067: d <= 8'h00;
                15'h4068: d <= 8'h00; 15'h4069: d <= 8'h00; 15'h406A: d <= 8'h00; 15'h406B: d <= 8'h00;
                15'h406C: d <= 8'h00; 15'h406D: d <= 8'h00; 15'h406E: d <= 8'h00; 15'h406F: d <= 8'h00;
                15'h4070: d <= 8'h00; 15'h4071: d <= 8'h00; 15'h4072: d <= 8'h00; 15'h4073: d <= 8'h00;
                15'h4074: d <= 8'h00; 15'h4075: d <= 8'h00; 15'h4076: d <= 8'h00; 15'h4077: d <= 8'h00;
                15'h4078: d <= 8'h00; 15'h4079: d <= 8'h00; 15'h407A: d <= 8'h00; 15'h407B: d <= 8'h00;
                15'h407C: d <= 8'h00; 15'h407D: d <= 8'h00; 15'h407E: d <= 8'h00; 15'h407F: d <= 8'hE0;
                15'h4080: d <= 8'h10; 15'h4081: d <= 8'h15; 15'h4082: d <= 8'h1A; 15'h4083: d <= 8'h1F;
                15'h4084: d <= 8'h20; 15'h4085: d <= 8'h25; 15'h4086: d <= 8'h2A; 15'h4087: d <= 8'h2F;
                15'h4088: d <= 8'h34; 15'h4089: d <= 8'h38; 15'h408A: d <= 8'h3C; 15'h408B: d <= 8'h31;
                15'h408C: d <= 8'h39; 15'h408D: d <= 8'h3D; 15'h408E: d <= 8'h32; 15'h408F: d <= 8'h36;
                15'h4090: d <= 8'h3E; 15'h4091: d <= 8'h33; 15'h4092: d <= 8'h37; 15'h4093: d <= 8'h3B;
                15'h4094: d <= 8'h44; 15'h4095: d <= 8'h48; 15'h4096: d <= 8'h4C; 15'h4097: d <= 8'h41;
                15'h4098: d <= 8'h49; 15'h4099: d <= 8'h4D; 15'h409A: d <= 8'h42; 15'h409B: d <= 8'h46;
                15'h409C: d <= 8'h4E; 15'h409D: d <= 8'h43; 15'h409E: d <= 8'h47; 15'h409F: d <= 8'h4B;
                15'h40A0: d <= 8'h50; 15'h40A1: d <= 8'h55; 15'h40A2: d <= 8'h5A; 15'h40A3: d <= 8'h5F;
                15'h40A4: d <= 8'h60; 15'h40A5: d <= 8'h65; 15'h40A6: d <= 8'h6A; 15'h40A7: d <= 8'h6F;
                15'h40A8: d <= 8'h74; 15'h40A9: d <= 8'h78; 15'h40AA: d <= 8'h7C; 15'h40AB: d <= 8'h71;
                15'h40AC: d <= 8'h79; 15'h40AD: d <= 8'h7D; 15'h40AE: d <= 8'h72; 15'h40AF: d <= 8'h76;
                15'h40B0: d <= 8'h7E; 15'h40B1: d <= 8'h73; 15'h40B2: d <= 8'h77; 15'h40B3: d <= 8'h7B;
                15'h40B4: d <= 8'h84; 15'h40B5: d <= 8'h88; 15'h40B6: d <= 8'h8C; 15'h40B7: d <= 8'h81;
                15'h40B8: d <= 8'h89; 15'h40B9: d <= 8'h8D; 15'h40BA: d <= 8'h82; 15'h40BB: d <= 8'h86;
                15'h40BC: d <= 8'h8E; 15'h40BD: d <= 8'h83; 15'h40BE: d <= 8'h87; 15'h40BF: d <= 8'h8B;
                15'h40C0: d <= 8'h90; 15'h40C1: d <= 8'h95; 15'h40C2: d <= 8'h9A; 15'h40C3: d <= 8'h9F;
                15'h40C4: d <= 8'hA4; 15'h40C5: d <= 8'hA8; 15'h40C6: d <= 8'hAC; 15'h40C7: d <= 8'hA1;
                15'h40C8: d <= 8'hA9; 15'h40C9: d <= 8'hAD; 15'h40CA: d <= 8'hA2; 15'h40CB: d <= 8'hA6;
                15'h40CC: d <= 8'hAE; 15'h40CD: d <= 8'hA3; 15'h40CE: d <= 8'hA7; 15'h40CF: d <= 8'hAB;
                15'h40D0: d <= 8'hB4; 15'h40D1: d <= 8'hB8; 15'h40D2: d <= 8'hBC; 15'h40D3: d <= 8'hB1;
                15'h40D4: d <= 8'hB9; 15'h40D5: d <= 8'hBD; 15'h40D6: d <= 8'hB2; 15'h40D7: d <= 8'hB6;
                15'h40D8: d <= 8'hBE; 15'h40D9: d <= 8'hB3; 15'h40DA: d <= 8'hB7; 15'h40DB: d <= 8'hBB;
                15'h40DC: d <= 8'hC4; 15'h40DD: d <= 8'hC8; 15'h40DE: d <= 8'hCC; 15'h40DF: d <= 8'hC1;
                15'h40E0: d <= 8'hC9; 15'h40E1: d <= 8'hCD; 15'h40E2: d <= 8'hC2; 15'h40E3: d <= 8'hC6;
                15'h40E4: d <= 8'hCE; 15'h40E5: d <= 8'hC3; 15'h40E6: d <= 8'hC7; 15'h40E7: d <= 8'hCB;
                15'h40E8: d <= 8'hC0; 15'h40E9: d <= 8'hC5; 15'h40EA: d <= 8'hCA; 15'h40EB: d <= 8'hCF;
                15'h40EC: d <= 8'hD0; 15'h40ED: d <= 8'hD5; 15'h40EE: d <= 8'hDA; 15'h40EF: d <= 8'hDF;
                15'h40F0: d <= 8'h74; 15'h40F1: d <= 8'h78; 15'h40F2: d <= 8'h7C; 15'h40F3: d <= 8'h71;
                15'h40F4: d <= 8'h79; 15'h40F5: d <= 8'h7D; 15'h40F6: d <= 8'h72; 15'h40F7: d <= 8'h76;
                15'h40F8: d <= 8'h7E; 15'h40F9: d <= 8'h73; 15'h40FA: d <= 8'h77; 15'h40FB: d <= 8'h7B;
                15'h40FC: d <= 8'hA0; 15'h40FD: d <= 8'hA5; 15'h40FE: d <= 8'hAA; 15'h40FF: d <= 8'hAF;
                15'h4100: d <= 8'h00; 15'h4101: d <= 8'h00; 15'h4102: d <= 8'h00; 15'h4103: d <= 8'h00;
                15'h4104: d <= 8'h00; 15'h4105: d <= 8'h00; 15'h4106: d <= 8'h00; 15'h4107: d <= 8'h00;
                15'h4108: d <= 8'h00; 15'h4109: d <= 8'h00; 15'h410A: d <= 8'h00; 15'h410B: d <= 8'h00;
                15'h410C: d <= 8'h00; 15'h410D: d <= 8'h00; 15'h410E: d <= 8'h00; 15'h410F: d <= 8'h00;
                15'h4110: d <= 8'h00; 15'h4111: d <= 8'h00; 15'h4112: d <= 8'h00; 15'h4113: d <= 8'h00;
                15'h4114: d <= 8'h00; 15'h4115: d <= 8'h00; 15'h4116: d <= 8'h00; 15'h4117: d <= 8'h00;
                15'h4118: d <= 8'h00; 15'h4119: d <= 8'h00; 15'h411A: d <= 8'h00; 15'h411B: d <= 8'h00;
                15'h411C: d <= 8'h00; 15'h411D: d <= 8'h00; 15'h411E: d <= 8'h00; 15'h411F: d <= 8'h00;
                15'h4120: d <= 8'h00; 15'h4121: d <= 8'h00; 15'h4122: d <= 8'h00; 15'h4123: d <= 8'h00;
                15'h4124: d <= 8'h00; 15'h4125: d <= 8'h00; 15'h4126: d <= 8'h00; 15'h4127: d <= 8'h00;
                15'h4128: d <= 8'h00; 15'h4129: d <= 8'h00; 15'h412A: d <= 8'h00; 15'h412B: d <= 8'h00;
                15'h412C: d <= 8'h00; 15'h412D: d <= 8'h00; 15'h412E: d <= 8'h00; 15'h412F: d <= 8'hAF;
                15'h4130: d <= 8'h00; 15'h4131: d <= 8'h00; 15'h4132: d <= 8'h00; 15'h4133: d <= 8'h00;
                15'h4134: d <= 8'h00; 15'h4135: d <= 8'h00; 15'h4136: d <= 8'h00; 15'h4137: d <= 8'h00;
                15'h4138: d <= 8'h00; 15'h4139: d <= 8'h00; 15'h413A: d <= 8'h00; 15'h413B: d <= 8'h00;
                15'h413C: d <= 8'h00; 15'h413D: d <= 8'h00; 15'h413E: d <= 8'h00; 15'h413F: d <= 8'h00;
                15'h4140: d <= 8'h00; 15'h4141: d <= 8'h00; 15'h4142: d <= 8'h00; 15'h4143: d <= 8'h00;
                15'h4144: d <= 8'h00; 15'h4145: d <= 8'h00; 15'h4146: d <= 8'h00; 15'h4147: d <= 8'h00;
                15'h4148: d <= 8'h00; 15'h4149: d <= 8'h00; 15'h414A: d <= 8'h00; 15'h414B: d <= 8'h00;
                15'h414C: d <= 8'h00; 15'h414D: d <= 8'h00; 15'h414E: d <= 8'h00; 15'h414F: d <= 8'h00;
                15'h4150: d <= 8'h00; 15'h4151: d <= 8'h00; 15'h4152: d <= 8'h00; 15'h4153: d <= 8'h00;
                15'h4154: d <= 8'h00; 15'h4155: d <= 8'h00; 15'h4156: d <= 8'h00; 15'h4157: d <= 8'h00;
                15'h4158: d <= 8'h45; 15'h4159: d <= 8'h35; 15'h415A: d <= 8'hAA; 15'h415B: d <= 8'h00;
                15'h415C: d <= 8'h00; 15'h415D: d <= 8'h00; 15'h415E: d <= 8'h00; 15'h415F: d <= 8'h00;
                15'h4160: d <= 8'h00; 15'h4161: d <= 8'h00; 15'h4162: d <= 8'h00; 15'h4163: d <= 8'h00;
                15'h4164: d <= 8'h00; 15'h4165: d <= 8'h00; 15'h4166: d <= 8'h00; 15'h4167: d <= 8'h00;
                15'h4168: d <= 8'h00; 15'h4169: d <= 8'h00; 15'h416A: d <= 8'h00; 15'h416B: d <= 8'h00;
                15'h416C: d <= 8'h00; 15'h416D: d <= 8'h00; 15'h416E: d <= 8'h00; 15'h416F: d <= 8'h00;
                15'h4170: d <= 8'h00; 15'h4171: d <= 8'h00; 15'h4172: d <= 8'h00; 15'h4173: d <= 8'h00;
                15'h4174: d <= 8'h00; 15'h4175: d <= 8'h00; 15'h4176: d <= 8'h00; 15'h4177: d <= 8'h00;
                15'h4178: d <= 8'h00; 15'h4179: d <= 8'h00; 15'h417A: d <= 8'h00; 15'h417B: d <= 8'h00;
                15'h417C: d <= 8'h00; 15'h417D: d <= 8'h00; 15'h417E: d <= 8'h00; 15'h417F: d <= 8'hE0;
                15'h4180: d <= 8'h10; 15'h4181: d <= 8'h15; 15'h4182: d <= 8'h1A; 15'h4183: d <= 8'h1F;
                15'h4184: d <= 8'h20; 15'h4185: d <= 8'h25; 15'h4186: d <= 8'h2A; 15'h4187: d <= 8'h2F;
                15'h4188: d <= 8'h34; 15'h4189: d <= 8'h38; 15'h418A: d <= 8'h3C; 15'h418B: d <= 8'h31;
                15'h418C: d <= 8'h39; 15'h418D: d <= 8'h3D; 15'h418E: d <= 8'h32; 15'h418F: d <= 8'h36;
                15'h4190: d <= 8'h3E; 15'h4191: d <= 8'h33; 15'h4192: d <= 8'h37; 15'h4193: d <= 8'h3B;
                15'h4194: d <= 8'h44; 15'h4195: d <= 8'h48; 15'h4196: d <= 8'h4C; 15'h4197: d <= 8'h41;
                15'h4198: d <= 8'h49; 15'h4199: d <= 8'h4D; 15'h419A: d <= 8'h42; 15'h419B: d <= 8'h46;
                15'h419C: d <= 8'h4E; 15'h419D: d <= 8'h43; 15'h419E: d <= 8'h47; 15'h419F: d <= 8'h4B;
                15'h41A0: d <= 8'h50; 15'h41A1: d <= 8'h55; 15'h41A2: d <= 8'h5A; 15'h41A3: d <= 8'h5F;
                15'h41A4: d <= 8'h60; 15'h41A5: d <= 8'h65; 15'h41A6: d <= 8'h6A; 15'h41A7: d <= 8'h6F;
                15'h41A8: d <= 8'h74; 15'h41A9: d <= 8'h78; 15'h41AA: d <= 8'h7C; 15'h41AB: d <= 8'h71;
                15'h41AC: d <= 8'h79; 15'h41AD: d <= 8'h7D; 15'h41AE: d <= 8'h72; 15'h41AF: d <= 8'h76;
                15'h41B0: d <= 8'h7E; 15'h41B1: d <= 8'h73; 15'h41B2: d <= 8'h77; 15'h41B3: d <= 8'h7B;
                15'h41B4: d <= 8'h84; 15'h41B5: d <= 8'h88; 15'h41B6: d <= 8'h8C; 15'h41B7: d <= 8'h81;
                15'h41B8: d <= 8'h89; 15'h41B9: d <= 8'h8D; 15'h41BA: d <= 8'h82; 15'h41BB: d <= 8'h86;
                15'h41BC: d <= 8'h8E; 15'h41BD: d <= 8'h83; 15'h41BE: d <= 8'h87; 15'h41BF: d <= 8'h8B;
                15'h41C0: d <= 8'h90; 15'h41C1: d <= 8'h95; 15'h41C2: d <= 8'h9A; 15'h41C3: d <= 8'h9F;
                15'h41C4: d <= 8'hA4; 15'h41C5: d <= 8'hA8; 15'h41C6: d <= 8'hAC; 15'h41C7: d <= 8'hA1;
                15'h41C8: d <= 8'hA9; 15'h41C9: d <= 8'hAD; 15'h41CA: d <= 8'hA2; 15'h41CB: d <= 8'hA6;
                15'h41CC: d <= 8'hAE; 15'h41CD: d <= 8'hA3; 15'h41CE: d <= 8'hA7; 15'h41CF: d <= 8'hAB;
                15'h41D0: d <= 8'hB4; 15'h41D1: d <= 8'hB8; 15'h41D2: d <= 8'hBC; 15'h41D3: d <= 8'hB1;
                15'h41D4: d <= 8'hB9; 15'h41D5: d <= 8'hBD; 15'h41D6: d <= 8'hB2; 15'h41D7: d <= 8'hB6;
                15'h41D8: d <= 8'hBE; 15'h41D9: d <= 8'hB3; 15'h41DA: d <= 8'hB7; 15'h41DB: d <= 8'hBB;
                15'h41DC: d <= 8'hC4; 15'h41DD: d <= 8'hC8; 15'h41DE: d <= 8'hCC; 15'h41DF: d <= 8'hC1;
                15'h41E0: d <= 8'hC9; 15'h41E1: d <= 8'hCD; 15'h41E2: d <= 8'hC2; 15'h41E3: d <= 8'hC6;
                15'h41E4: d <= 8'hCE; 15'h41E5: d <= 8'hC3; 15'h41E6: d <= 8'hC7; 15'h41E7: d <= 8'hCB;
                15'h41E8: d <= 8'hC0; 15'h41E9: d <= 8'hC5; 15'h41EA: d <= 8'hCA; 15'h41EB: d <= 8'hCF;
                15'h41EC: d <= 8'hD0; 15'h41ED: d <= 8'hD5; 15'h41EE: d <= 8'hDA; 15'h41EF: d <= 8'hDF;
                15'h41F0: d <= 8'h74; 15'h41F1: d <= 8'h78; 15'h41F2: d <= 8'h7C; 15'h41F3: d <= 8'h71;
                15'h41F4: d <= 8'h79; 15'h41F5: d <= 8'h7D; 15'h41F6: d <= 8'h72; 15'h41F7: d <= 8'h76;
                15'h41F8: d <= 8'h7E; 15'h41F9: d <= 8'h73; 15'h41FA: d <= 8'h77; 15'h41FB: d <= 8'h7B;
                15'h41FC: d <= 8'hA0; 15'h41FD: d <= 8'hA5; 15'h41FE: d <= 8'hAA; 15'h41FF: d <= 8'hAF;
                15'h4200: d <= 8'h00; 15'h4201: d <= 8'h00; 15'h4202: d <= 8'h00; 15'h4203: d <= 8'h00;
                15'h4204: d <= 8'h00; 15'h4205: d <= 8'h00; 15'h4206: d <= 8'h00; 15'h4207: d <= 8'h00;
                15'h4208: d <= 8'h00; 15'h4209: d <= 8'h00; 15'h420A: d <= 8'h00; 15'h420B: d <= 8'h00;
                15'h420C: d <= 8'h00; 15'h420D: d <= 8'h00; 15'h420E: d <= 8'h00; 15'h420F: d <= 8'h00;
                15'h4210: d <= 8'h00; 15'h4211: d <= 8'h00; 15'h4212: d <= 8'h00; 15'h4213: d <= 8'h00;
                15'h4214: d <= 8'h00; 15'h4215: d <= 8'h00; 15'h4216: d <= 8'h00; 15'h4217: d <= 8'h00;
                15'h4218: d <= 8'h00; 15'h4219: d <= 8'h00; 15'h421A: d <= 8'h00; 15'h421B: d <= 8'h00;
                15'h421C: d <= 8'h00; 15'h421D: d <= 8'h00; 15'h421E: d <= 8'h00; 15'h421F: d <= 8'h00;
                15'h4220: d <= 8'h00; 15'h4221: d <= 8'h00; 15'h4222: d <= 8'h00; 15'h4223: d <= 8'h00;
                15'h4224: d <= 8'h00; 15'h4225: d <= 8'h00; 15'h4226: d <= 8'h00; 15'h4227: d <= 8'h00;
                15'h4228: d <= 8'h00; 15'h4229: d <= 8'h00; 15'h422A: d <= 8'h00; 15'h422B: d <= 8'h00;
                15'h422C: d <= 8'h00; 15'h422D: d <= 8'h00; 15'h422E: d <= 8'h00; 15'h422F: d <= 8'hAF;
                15'h4230: d <= 8'h00; 15'h4231: d <= 8'h00; 15'h4232: d <= 8'h00; 15'h4233: d <= 8'h00;
                15'h4234: d <= 8'h00; 15'h4235: d <= 8'h00; 15'h4236: d <= 8'h00; 15'h4237: d <= 8'h00;
                15'h4238: d <= 8'h00; 15'h4239: d <= 8'h00; 15'h423A: d <= 8'h00; 15'h423B: d <= 8'h00;
                15'h423C: d <= 8'h00; 15'h423D: d <= 8'h00; 15'h423E: d <= 8'h00; 15'h423F: d <= 8'h00;
                15'h4240: d <= 8'h00; 15'h4241: d <= 8'h00; 15'h4242: d <= 8'h00; 15'h4243: d <= 8'h00;
                15'h4244: d <= 8'h00; 15'h4245: d <= 8'h00; 15'h4246: d <= 8'h00; 15'h4247: d <= 8'h00;
                15'h4248: d <= 8'h00; 15'h4249: d <= 8'h00; 15'h424A: d <= 8'h00; 15'h424B: d <= 8'h00;
                15'h424C: d <= 8'h00; 15'h424D: d <= 8'h00; 15'h424E: d <= 8'h00; 15'h424F: d <= 8'h00;
                15'h4250: d <= 8'h00; 15'h4251: d <= 8'h00; 15'h4252: d <= 8'h00; 15'h4253: d <= 8'h00;
                15'h4254: d <= 8'h00; 15'h4255: d <= 8'h00; 15'h4256: d <= 8'h00; 15'h4257: d <= 8'h00;
                15'h4258: d <= 8'h45; 15'h4259: d <= 8'h35; 15'h425A: d <= 8'hAA; 15'h425B: d <= 8'h00;
                15'h425C: d <= 8'h00; 15'h425D: d <= 8'h00; 15'h425E: d <= 8'h00; 15'h425F: d <= 8'h00;
                15'h4260: d <= 8'h00; 15'h4261: d <= 8'h00; 15'h4262: d <= 8'h00; 15'h4263: d <= 8'h00;
                15'h4264: d <= 8'h00; 15'h4265: d <= 8'h00; 15'h4266: d <= 8'h00; 15'h4267: d <= 8'h00;
                15'h4268: d <= 8'h00; 15'h4269: d <= 8'h00; 15'h426A: d <= 8'h00; 15'h426B: d <= 8'h00;
                15'h426C: d <= 8'h00; 15'h426D: d <= 8'h00; 15'h426E: d <= 8'h00; 15'h426F: d <= 8'h00;
                15'h4270: d <= 8'h00; 15'h4271: d <= 8'h00; 15'h4272: d <= 8'h00; 15'h4273: d <= 8'h00;
                15'h4274: d <= 8'h00; 15'h4275: d <= 8'h00; 15'h4276: d <= 8'h00; 15'h4277: d <= 8'h00;
                15'h4278: d <= 8'h00; 15'h4279: d <= 8'h00; 15'h427A: d <= 8'h00; 15'h427B: d <= 8'h00;
                15'h427C: d <= 8'h00; 15'h427D: d <= 8'h00; 15'h427E: d <= 8'h00; 15'h427F: d <= 8'hE0;
                15'h4280: d <= 8'h10; 15'h4281: d <= 8'h15; 15'h4282: d <= 8'h1A; 15'h4283: d <= 8'h1F;
                15'h4284: d <= 8'h20; 15'h4285: d <= 8'h25; 15'h4286: d <= 8'h2A; 15'h4287: d <= 8'h2F;
                15'h4288: d <= 8'h34; 15'h4289: d <= 8'h38; 15'h428A: d <= 8'h3C; 15'h428B: d <= 8'h31;
                15'h428C: d <= 8'h39; 15'h428D: d <= 8'h3D; 15'h428E: d <= 8'h32; 15'h428F: d <= 8'h36;
                15'h4290: d <= 8'h3E; 15'h4291: d <= 8'h33; 15'h4292: d <= 8'h37; 15'h4293: d <= 8'h3B;
                15'h4294: d <= 8'h44; 15'h4295: d <= 8'h48; 15'h4296: d <= 8'h4C; 15'h4297: d <= 8'h41;
                15'h4298: d <= 8'h49; 15'h4299: d <= 8'h4D; 15'h429A: d <= 8'h42; 15'h429B: d <= 8'h46;
                15'h429C: d <= 8'h4E; 15'h429D: d <= 8'h43; 15'h429E: d <= 8'h47; 15'h429F: d <= 8'h4B;
                15'h42A0: d <= 8'h50; 15'h42A1: d <= 8'h55; 15'h42A2: d <= 8'h5A; 15'h42A3: d <= 8'h5F;
                15'h42A4: d <= 8'h60; 15'h42A5: d <= 8'h65; 15'h42A6: d <= 8'h6A; 15'h42A7: d <= 8'h6F;
                15'h42A8: d <= 8'h74; 15'h42A9: d <= 8'h78; 15'h42AA: d <= 8'h7C; 15'h42AB: d <= 8'h71;
                15'h42AC: d <= 8'h79; 15'h42AD: d <= 8'h7D; 15'h42AE: d <= 8'h72; 15'h42AF: d <= 8'h76;
                15'h42B0: d <= 8'h7E; 15'h42B1: d <= 8'h73; 15'h42B2: d <= 8'h77; 15'h42B3: d <= 8'h7B;
                15'h42B4: d <= 8'h84; 15'h42B5: d <= 8'h88; 15'h42B6: d <= 8'h8C; 15'h42B7: d <= 8'h81;
                15'h42B8: d <= 8'h89; 15'h42B9: d <= 8'h8D; 15'h42BA: d <= 8'h82; 15'h42BB: d <= 8'h86;
                15'h42BC: d <= 8'h8E; 15'h42BD: d <= 8'h83; 15'h42BE: d <= 8'h87; 15'h42BF: d <= 8'h8B;
                15'h42C0: d <= 8'h90; 15'h42C1: d <= 8'h95; 15'h42C2: d <= 8'h9A; 15'h42C3: d <= 8'h9F;
                15'h42C4: d <= 8'hA4; 15'h42C5: d <= 8'hA8; 15'h42C6: d <= 8'hAC; 15'h42C7: d <= 8'hA1;
                15'h42C8: d <= 8'hA9; 15'h42C9: d <= 8'hAD; 15'h42CA: d <= 8'hA2; 15'h42CB: d <= 8'hA6;
                15'h42CC: d <= 8'hAE; 15'h42CD: d <= 8'hA3; 15'h42CE: d <= 8'hA7; 15'h42CF: d <= 8'hAB;
                15'h42D0: d <= 8'hB4; 15'h42D1: d <= 8'hB8; 15'h42D2: d <= 8'hBC; 15'h42D3: d <= 8'hB1;
                15'h42D4: d <= 8'hB9; 15'h42D5: d <= 8'hBD; 15'h42D6: d <= 8'hB2; 15'h42D7: d <= 8'hB6;
                15'h42D8: d <= 8'hBE; 15'h42D9: d <= 8'hB3; 15'h42DA: d <= 8'hB7; 15'h42DB: d <= 8'hBB;
                15'h42DC: d <= 8'hC4; 15'h42DD: d <= 8'hC8; 15'h42DE: d <= 8'hCC; 15'h42DF: d <= 8'hC1;
                15'h42E0: d <= 8'hC9; 15'h42E1: d <= 8'hCD; 15'h42E2: d <= 8'hC2; 15'h42E3: d <= 8'hC6;
                15'h42E4: d <= 8'hCE; 15'h42E5: d <= 8'hC3; 15'h42E6: d <= 8'hC7; 15'h42E7: d <= 8'hCB;
                15'h42E8: d <= 8'hC0; 15'h42E9: d <= 8'hC5; 15'h42EA: d <= 8'hCA; 15'h42EB: d <= 8'hCF;
                15'h42EC: d <= 8'hD0; 15'h42ED: d <= 8'hD5; 15'h42EE: d <= 8'hDA; 15'h42EF: d <= 8'hDF;
                15'h42F0: d <= 8'h74; 15'h42F1: d <= 8'h78; 15'h42F2: d <= 8'h7C; 15'h42F3: d <= 8'h71;
                15'h42F4: d <= 8'h79; 15'h42F5: d <= 8'h7D; 15'h42F6: d <= 8'h72; 15'h42F7: d <= 8'h76;
                15'h42F8: d <= 8'h7E; 15'h42F9: d <= 8'h73; 15'h42FA: d <= 8'h77; 15'h42FB: d <= 8'h7B;
                15'h42FC: d <= 8'hA0; 15'h42FD: d <= 8'hA5; 15'h42FE: d <= 8'hAA; 15'h42FF: d <= 8'hAF;
                15'h4300: d <= 8'h00; 15'h4301: d <= 8'h00; 15'h4302: d <= 8'h00; 15'h4303: d <= 8'h00;
                15'h4304: d <= 8'h00; 15'h4305: d <= 8'h00; 15'h4306: d <= 8'h00; 15'h4307: d <= 8'h00;
                15'h4308: d <= 8'h00; 15'h4309: d <= 8'h00; 15'h430A: d <= 8'h00; 15'h430B: d <= 8'h00;
                15'h430C: d <= 8'h00; 15'h430D: d <= 8'h00; 15'h430E: d <= 8'h00; 15'h430F: d <= 8'h00;
                15'h4310: d <= 8'h00; 15'h4311: d <= 8'h00; 15'h4312: d <= 8'h00; 15'h4313: d <= 8'h00;
                15'h4314: d <= 8'h00; 15'h4315: d <= 8'h00; 15'h4316: d <= 8'h00; 15'h4317: d <= 8'h00;
                15'h4318: d <= 8'h00; 15'h4319: d <= 8'h00; 15'h431A: d <= 8'h00; 15'h431B: d <= 8'h00;
                15'h431C: d <= 8'h00; 15'h431D: d <= 8'h00; 15'h431E: d <= 8'h00; 15'h431F: d <= 8'h00;
                15'h4320: d <= 8'h00; 15'h4321: d <= 8'h00; 15'h4322: d <= 8'h00; 15'h4323: d <= 8'h00;
                15'h4324: d <= 8'h00; 15'h4325: d <= 8'h00; 15'h4326: d <= 8'h00; 15'h4327: d <= 8'h00;
                15'h4328: d <= 8'h00; 15'h4329: d <= 8'h00; 15'h432A: d <= 8'h00; 15'h432B: d <= 8'h00;
                15'h432C: d <= 8'h00; 15'h432D: d <= 8'h00; 15'h432E: d <= 8'h00; 15'h432F: d <= 8'hAF;
                15'h4330: d <= 8'h00; 15'h4331: d <= 8'h00; 15'h4332: d <= 8'h00; 15'h4333: d <= 8'h00;
                15'h4334: d <= 8'h00; 15'h4335: d <= 8'h00; 15'h4336: d <= 8'h00; 15'h4337: d <= 8'h00;
                15'h4338: d <= 8'h00; 15'h4339: d <= 8'h00; 15'h433A: d <= 8'h00; 15'h433B: d <= 8'h00;
                15'h433C: d <= 8'h00; 15'h433D: d <= 8'h00; 15'h433E: d <= 8'h00; 15'h433F: d <= 8'h00;
                15'h4340: d <= 8'h00; 15'h4341: d <= 8'h00; 15'h4342: d <= 8'h00; 15'h4343: d <= 8'h00;
                15'h4344: d <= 8'h00; 15'h4345: d <= 8'h00; 15'h4346: d <= 8'h00; 15'h4347: d <= 8'h00;
                15'h4348: d <= 8'h00; 15'h4349: d <= 8'h00; 15'h434A: d <= 8'h00; 15'h434B: d <= 8'h00;
                15'h434C: d <= 8'h00; 15'h434D: d <= 8'h00; 15'h434E: d <= 8'h00; 15'h434F: d <= 8'h00;
                15'h4350: d <= 8'h00; 15'h4351: d <= 8'h00; 15'h4352: d <= 8'h00; 15'h4353: d <= 8'h00;
                15'h4354: d <= 8'h00; 15'h4355: d <= 8'h00; 15'h4356: d <= 8'h00; 15'h4357: d <= 8'h00;
                15'h4358: d <= 8'h45; 15'h4359: d <= 8'h35; 15'h435A: d <= 8'hAA; 15'h435B: d <= 8'h00;
                15'h435C: d <= 8'h00; 15'h435D: d <= 8'h00; 15'h435E: d <= 8'h00; 15'h435F: d <= 8'h00;
                15'h4360: d <= 8'h00; 15'h4361: d <= 8'h00; 15'h4362: d <= 8'h00; 15'h4363: d <= 8'h00;
                15'h4364: d <= 8'h00; 15'h4365: d <= 8'h00; 15'h4366: d <= 8'h00; 15'h4367: d <= 8'h00;
                15'h4368: d <= 8'h00; 15'h4369: d <= 8'h00; 15'h436A: d <= 8'h00; 15'h436B: d <= 8'h00;
                15'h436C: d <= 8'h00; 15'h436D: d <= 8'h00; 15'h436E: d <= 8'h00; 15'h436F: d <= 8'h00;
                15'h4370: d <= 8'h00; 15'h4371: d <= 8'h00; 15'h4372: d <= 8'h00; 15'h4373: d <= 8'h00;
                15'h4374: d <= 8'h00; 15'h4375: d <= 8'h00; 15'h4376: d <= 8'h00; 15'h4377: d <= 8'h00;
                15'h4378: d <= 8'h00; 15'h4379: d <= 8'h00; 15'h437A: d <= 8'h00; 15'h437B: d <= 8'h00;
                15'h437C: d <= 8'h00; 15'h437D: d <= 8'h00; 15'h437E: d <= 8'h00; 15'h437F: d <= 8'hE0;
                15'h4380: d <= 8'h10; 15'h4381: d <= 8'h15; 15'h4382: d <= 8'h1A; 15'h4383: d <= 8'h1F;
                15'h4384: d <= 8'h20; 15'h4385: d <= 8'h25; 15'h4386: d <= 8'h2A; 15'h4387: d <= 8'h2F;
                15'h4388: d <= 8'h34; 15'h4389: d <= 8'h38; 15'h438A: d <= 8'h3C; 15'h438B: d <= 8'h31;
                15'h438C: d <= 8'h39; 15'h438D: d <= 8'h3D; 15'h438E: d <= 8'h32; 15'h438F: d <= 8'h36;
                15'h4390: d <= 8'h3E; 15'h4391: d <= 8'h33; 15'h4392: d <= 8'h37; 15'h4393: d <= 8'h3B;
                15'h4394: d <= 8'h44; 15'h4395: d <= 8'h48; 15'h4396: d <= 8'h4C; 15'h4397: d <= 8'h41;
                15'h4398: d <= 8'h49; 15'h4399: d <= 8'h4D; 15'h439A: d <= 8'h42; 15'h439B: d <= 8'h46;
                15'h439C: d <= 8'h4E; 15'h439D: d <= 8'h43; 15'h439E: d <= 8'h47; 15'h439F: d <= 8'h4B;
                15'h43A0: d <= 8'h50; 15'h43A1: d <= 8'h55; 15'h43A2: d <= 8'h5A; 15'h43A3: d <= 8'h5F;
                15'h43A4: d <= 8'h60; 15'h43A5: d <= 8'h65; 15'h43A6: d <= 8'h6A; 15'h43A7: d <= 8'h6F;
                15'h43A8: d <= 8'h74; 15'h43A9: d <= 8'h78; 15'h43AA: d <= 8'h7C; 15'h43AB: d <= 8'h71;
                15'h43AC: d <= 8'h79; 15'h43AD: d <= 8'h7D; 15'h43AE: d <= 8'h72; 15'h43AF: d <= 8'h76;
                15'h43B0: d <= 8'h7E; 15'h43B1: d <= 8'h73; 15'h43B2: d <= 8'h77; 15'h43B3: d <= 8'h7B;
                15'h43B4: d <= 8'h84; 15'h43B5: d <= 8'h88; 15'h43B6: d <= 8'h8C; 15'h43B7: d <= 8'h81;
                15'h43B8: d <= 8'h89; 15'h43B9: d <= 8'h8D; 15'h43BA: d <= 8'h82; 15'h43BB: d <= 8'h86;
                15'h43BC: d <= 8'h8E; 15'h43BD: d <= 8'h83; 15'h43BE: d <= 8'h87; 15'h43BF: d <= 8'h8B;
                15'h43C0: d <= 8'h90; 15'h43C1: d <= 8'h95; 15'h43C2: d <= 8'h9A; 15'h43C3: d <= 8'h9F;
                15'h43C4: d <= 8'hA4; 15'h43C5: d <= 8'hA8; 15'h43C6: d <= 8'hAC; 15'h43C7: d <= 8'hA1;
                15'h43C8: d <= 8'hA9; 15'h43C9: d <= 8'hAD; 15'h43CA: d <= 8'hA2; 15'h43CB: d <= 8'hA6;
                15'h43CC: d <= 8'hAE; 15'h43CD: d <= 8'hA3; 15'h43CE: d <= 8'hA7; 15'h43CF: d <= 8'hAB;
                15'h43D0: d <= 8'hB4; 15'h43D1: d <= 8'hB8; 15'h43D2: d <= 8'hBC; 15'h43D3: d <= 8'hB1;
                15'h43D4: d <= 8'hB9; 15'h43D5: d <= 8'hBD; 15'h43D6: d <= 8'hB2; 15'h43D7: d <= 8'hB6;
                15'h43D8: d <= 8'hBE; 15'h43D9: d <= 8'hB3; 15'h43DA: d <= 8'hB7; 15'h43DB: d <= 8'hBB;
                15'h43DC: d <= 8'hC4; 15'h43DD: d <= 8'hC8; 15'h43DE: d <= 8'hCC; 15'h43DF: d <= 8'hC1;
                15'h43E0: d <= 8'hC9; 15'h43E1: d <= 8'hCD; 15'h43E2: d <= 8'hC2; 15'h43E3: d <= 8'hC6;
                15'h43E4: d <= 8'hCE; 15'h43E5: d <= 8'hC3; 15'h43E6: d <= 8'hC7; 15'h43E7: d <= 8'hCB;
                15'h43E8: d <= 8'hC0; 15'h43E9: d <= 8'hC5; 15'h43EA: d <= 8'hCA; 15'h43EB: d <= 8'hCF;
                15'h43EC: d <= 8'hD0; 15'h43ED: d <= 8'hD5; 15'h43EE: d <= 8'hDA; 15'h43EF: d <= 8'hDF;
                15'h43F0: d <= 8'h74; 15'h43F1: d <= 8'h78; 15'h43F2: d <= 8'h7C; 15'h43F3: d <= 8'h71;
                15'h43F4: d <= 8'h79; 15'h43F5: d <= 8'h7D; 15'h43F6: d <= 8'h72; 15'h43F7: d <= 8'h76;
                15'h43F8: d <= 8'h7E; 15'h43F9: d <= 8'h73; 15'h43FA: d <= 8'h77; 15'h43FB: d <= 8'h7B;
                15'h43FC: d <= 8'hA0; 15'h43FD: d <= 8'hA5; 15'h43FE: d <= 8'hAA; 15'h43FF: d <= 8'hAF;
                15'h4400: d <= 8'h00; 15'h4401: d <= 8'h00; 15'h4402: d <= 8'h00; 15'h4403: d <= 8'h00;
                15'h4404: d <= 8'h00; 15'h4405: d <= 8'h00; 15'h4406: d <= 8'h00; 15'h4407: d <= 8'h00;
                15'h4408: d <= 8'h00; 15'h4409: d <= 8'h00; 15'h440A: d <= 8'h00; 15'h440B: d <= 8'h00;
                15'h440C: d <= 8'h00; 15'h440D: d <= 8'h00; 15'h440E: d <= 8'h00; 15'h440F: d <= 8'h00;
                15'h4410: d <= 8'h00; 15'h4411: d <= 8'h00; 15'h4412: d <= 8'h00; 15'h4413: d <= 8'h00;
                15'h4414: d <= 8'h00; 15'h4415: d <= 8'h00; 15'h4416: d <= 8'h00; 15'h4417: d <= 8'h00;
                15'h4418: d <= 8'h00; 15'h4419: d <= 8'h00; 15'h441A: d <= 8'h00; 15'h441B: d <= 8'h00;
                15'h441C: d <= 8'h00; 15'h441D: d <= 8'h00; 15'h441E: d <= 8'h00; 15'h441F: d <= 8'h00;
                15'h4420: d <= 8'h00; 15'h4421: d <= 8'h00; 15'h4422: d <= 8'h00; 15'h4423: d <= 8'h00;
                15'h4424: d <= 8'h00; 15'h4425: d <= 8'h00; 15'h4426: d <= 8'h00; 15'h4427: d <= 8'h00;
                15'h4428: d <= 8'h00; 15'h4429: d <= 8'h00; 15'h442A: d <= 8'h00; 15'h442B: d <= 8'h00;
                15'h442C: d <= 8'h00; 15'h442D: d <= 8'h00; 15'h442E: d <= 8'h00; 15'h442F: d <= 8'hAF;
                15'h4430: d <= 8'h00; 15'h4431: d <= 8'h00; 15'h4432: d <= 8'h00; 15'h4433: d <= 8'h00;
                15'h4434: d <= 8'h00; 15'h4435: d <= 8'h00; 15'h4436: d <= 8'h00; 15'h4437: d <= 8'h00;
                15'h4438: d <= 8'h00; 15'h4439: d <= 8'h00; 15'h443A: d <= 8'h00; 15'h443B: d <= 8'h00;
                15'h443C: d <= 8'h00; 15'h443D: d <= 8'h00; 15'h443E: d <= 8'h00; 15'h443F: d <= 8'h00;
                15'h4440: d <= 8'h00; 15'h4441: d <= 8'h00; 15'h4442: d <= 8'h00; 15'h4443: d <= 8'h00;
                15'h4444: d <= 8'h00; 15'h4445: d <= 8'h00; 15'h4446: d <= 8'h00; 15'h4447: d <= 8'h00;
                15'h4448: d <= 8'h00; 15'h4449: d <= 8'h00; 15'h444A: d <= 8'h00; 15'h444B: d <= 8'h00;
                15'h444C: d <= 8'h00; 15'h444D: d <= 8'h00; 15'h444E: d <= 8'h00; 15'h444F: d <= 8'h00;
                15'h4450: d <= 8'h00; 15'h4451: d <= 8'h00; 15'h4452: d <= 8'h00; 15'h4453: d <= 8'h00;
                15'h4454: d <= 8'h00; 15'h4455: d <= 8'h00; 15'h4456: d <= 8'h00; 15'h4457: d <= 8'h00;
                15'h4458: d <= 8'h45; 15'h4459: d <= 8'h35; 15'h445A: d <= 8'hAA; 15'h445B: d <= 8'h00;
                15'h445C: d <= 8'h00; 15'h445D: d <= 8'h00; 15'h445E: d <= 8'h00; 15'h445F: d <= 8'h00;
                15'h4460: d <= 8'h00; 15'h4461: d <= 8'h00; 15'h4462: d <= 8'h00; 15'h4463: d <= 8'h00;
                15'h4464: d <= 8'h00; 15'h4465: d <= 8'h00; 15'h4466: d <= 8'h00; 15'h4467: d <= 8'h00;
                15'h4468: d <= 8'h00; 15'h4469: d <= 8'h00; 15'h446A: d <= 8'h00; 15'h446B: d <= 8'h00;
                15'h446C: d <= 8'h00; 15'h446D: d <= 8'h00; 15'h446E: d <= 8'h00; 15'h446F: d <= 8'h00;
                15'h4470: d <= 8'h00; 15'h4471: d <= 8'h00; 15'h4472: d <= 8'h00; 15'h4473: d <= 8'h00;
                15'h4474: d <= 8'h00; 15'h4475: d <= 8'h00; 15'h4476: d <= 8'h00; 15'h4477: d <= 8'h00;
                15'h4478: d <= 8'h00; 15'h4479: d <= 8'h00; 15'h447A: d <= 8'h00; 15'h447B: d <= 8'h00;
                15'h447C: d <= 8'h00; 15'h447D: d <= 8'h00; 15'h447E: d <= 8'h00; 15'h447F: d <= 8'hE0;
                15'h4480: d <= 8'h10; 15'h4481: d <= 8'h15; 15'h4482: d <= 8'h1A; 15'h4483: d <= 8'h1F;
                15'h4484: d <= 8'h20; 15'h4485: d <= 8'h25; 15'h4486: d <= 8'h2A; 15'h4487: d <= 8'h2F;
                15'h4488: d <= 8'h34; 15'h4489: d <= 8'h38; 15'h448A: d <= 8'h3C; 15'h448B: d <= 8'h31;
                15'h448C: d <= 8'h39; 15'h448D: d <= 8'h3D; 15'h448E: d <= 8'h32; 15'h448F: d <= 8'h36;
                15'h4490: d <= 8'h3E; 15'h4491: d <= 8'h33; 15'h4492: d <= 8'h37; 15'h4493: d <= 8'h3B;
                15'h4494: d <= 8'h44; 15'h4495: d <= 8'h48; 15'h4496: d <= 8'h4C; 15'h4497: d <= 8'h41;
                15'h4498: d <= 8'h49; 15'h4499: d <= 8'h4D; 15'h449A: d <= 8'h42; 15'h449B: d <= 8'h46;
                15'h449C: d <= 8'h4E; 15'h449D: d <= 8'h43; 15'h449E: d <= 8'h47; 15'h449F: d <= 8'h4B;
                15'h44A0: d <= 8'h50; 15'h44A1: d <= 8'h55; 15'h44A2: d <= 8'h5A; 15'h44A3: d <= 8'h5F;
                15'h44A4: d <= 8'h60; 15'h44A5: d <= 8'h65; 15'h44A6: d <= 8'h6A; 15'h44A7: d <= 8'h6F;
                15'h44A8: d <= 8'h74; 15'h44A9: d <= 8'h78; 15'h44AA: d <= 8'h7C; 15'h44AB: d <= 8'h71;
                15'h44AC: d <= 8'h79; 15'h44AD: d <= 8'h7D; 15'h44AE: d <= 8'h72; 15'h44AF: d <= 8'h76;
                15'h44B0: d <= 8'h7E; 15'h44B1: d <= 8'h73; 15'h44B2: d <= 8'h77; 15'h44B3: d <= 8'h7B;
                15'h44B4: d <= 8'h84; 15'h44B5: d <= 8'h88; 15'h44B6: d <= 8'h8C; 15'h44B7: d <= 8'h81;
                15'h44B8: d <= 8'h89; 15'h44B9: d <= 8'h8D; 15'h44BA: d <= 8'h82; 15'h44BB: d <= 8'h86;
                15'h44BC: d <= 8'h8E; 15'h44BD: d <= 8'h83; 15'h44BE: d <= 8'h87; 15'h44BF: d <= 8'h8B;
                15'h44C0: d <= 8'h90; 15'h44C1: d <= 8'h95; 15'h44C2: d <= 8'h9A; 15'h44C3: d <= 8'h9F;
                15'h44C4: d <= 8'hA4; 15'h44C5: d <= 8'hA8; 15'h44C6: d <= 8'hAC; 15'h44C7: d <= 8'hA1;
                15'h44C8: d <= 8'hA9; 15'h44C9: d <= 8'hAD; 15'h44CA: d <= 8'hA2; 15'h44CB: d <= 8'hA6;
                15'h44CC: d <= 8'hAE; 15'h44CD: d <= 8'hA3; 15'h44CE: d <= 8'hA7; 15'h44CF: d <= 8'hAB;
                15'h44D0: d <= 8'hB4; 15'h44D1: d <= 8'hB8; 15'h44D2: d <= 8'hBC; 15'h44D3: d <= 8'hB1;
                15'h44D4: d <= 8'hB9; 15'h44D5: d <= 8'hBD; 15'h44D6: d <= 8'hB2; 15'h44D7: d <= 8'hB6;
                15'h44D8: d <= 8'hBE; 15'h44D9: d <= 8'hB3; 15'h44DA: d <= 8'hB7; 15'h44DB: d <= 8'hBB;
                15'h44DC: d <= 8'hC4; 15'h44DD: d <= 8'hC8; 15'h44DE: d <= 8'hCC; 15'h44DF: d <= 8'hC1;
                15'h44E0: d <= 8'hC9; 15'h44E1: d <= 8'hCD; 15'h44E2: d <= 8'hC2; 15'h44E3: d <= 8'hC6;
                15'h44E4: d <= 8'hCE; 15'h44E5: d <= 8'hC3; 15'h44E6: d <= 8'hC7; 15'h44E7: d <= 8'hCB;
                15'h44E8: d <= 8'hC0; 15'h44E9: d <= 8'hC5; 15'h44EA: d <= 8'hCA; 15'h44EB: d <= 8'hCF;
                15'h44EC: d <= 8'hD0; 15'h44ED: d <= 8'hD5; 15'h44EE: d <= 8'hDA; 15'h44EF: d <= 8'hDF;
                15'h44F0: d <= 8'h74; 15'h44F1: d <= 8'h78; 15'h44F2: d <= 8'h7C; 15'h44F3: d <= 8'h71;
                15'h44F4: d <= 8'h79; 15'h44F5: d <= 8'h7D; 15'h44F6: d <= 8'h72; 15'h44F7: d <= 8'h76;
                15'h44F8: d <= 8'h7E; 15'h44F9: d <= 8'h73; 15'h44FA: d <= 8'h77; 15'h44FB: d <= 8'h7B;
                15'h44FC: d <= 8'hA0; 15'h44FD: d <= 8'hA5; 15'h44FE: d <= 8'hAA; 15'h44FF: d <= 8'hAF;
                15'h4500: d <= 8'h00; 15'h4501: d <= 8'h00; 15'h4502: d <= 8'h00; 15'h4503: d <= 8'h00;
                15'h4504: d <= 8'h00; 15'h4505: d <= 8'h00; 15'h4506: d <= 8'h00; 15'h4507: d <= 8'h00;
                15'h4508: d <= 8'h00; 15'h4509: d <= 8'h00; 15'h450A: d <= 8'h00; 15'h450B: d <= 8'h00;
                15'h450C: d <= 8'h00; 15'h450D: d <= 8'h00; 15'h450E: d <= 8'h00; 15'h450F: d <= 8'h00;
                15'h4510: d <= 8'h00; 15'h4511: d <= 8'h00; 15'h4512: d <= 8'h00; 15'h4513: d <= 8'h00;
                15'h4514: d <= 8'h00; 15'h4515: d <= 8'h00; 15'h4516: d <= 8'h00; 15'h4517: d <= 8'h00;
                15'h4518: d <= 8'h00; 15'h4519: d <= 8'h00; 15'h451A: d <= 8'h00; 15'h451B: d <= 8'h00;
                15'h451C: d <= 8'h00; 15'h451D: d <= 8'h00; 15'h451E: d <= 8'h00; 15'h451F: d <= 8'h00;
                15'h4520: d <= 8'h00; 15'h4521: d <= 8'h00; 15'h4522: d <= 8'h00; 15'h4523: d <= 8'h00;
                15'h4524: d <= 8'h00; 15'h4525: d <= 8'h00; 15'h4526: d <= 8'h00; 15'h4527: d <= 8'h00;
                15'h4528: d <= 8'h00; 15'h4529: d <= 8'h00; 15'h452A: d <= 8'h00; 15'h452B: d <= 8'h00;
                15'h452C: d <= 8'h00; 15'h452D: d <= 8'h00; 15'h452E: d <= 8'h00; 15'h452F: d <= 8'hAF;
                15'h4530: d <= 8'h00; 15'h4531: d <= 8'h00; 15'h4532: d <= 8'h00; 15'h4533: d <= 8'h00;
                15'h4534: d <= 8'h00; 15'h4535: d <= 8'h00; 15'h4536: d <= 8'h00; 15'h4537: d <= 8'h00;
                15'h4538: d <= 8'h00; 15'h4539: d <= 8'h00; 15'h453A: d <= 8'h00; 15'h453B: d <= 8'h00;
                15'h453C: d <= 8'h00; 15'h453D: d <= 8'h00; 15'h453E: d <= 8'h00; 15'h453F: d <= 8'h00;
                15'h4540: d <= 8'h00; 15'h4541: d <= 8'h00; 15'h4542: d <= 8'h00; 15'h4543: d <= 8'h00;
                15'h4544: d <= 8'h00; 15'h4545: d <= 8'h00; 15'h4546: d <= 8'h00; 15'h4547: d <= 8'h00;
                15'h4548: d <= 8'h00; 15'h4549: d <= 8'h00; 15'h454A: d <= 8'h00; 15'h454B: d <= 8'h00;
                15'h454C: d <= 8'h00; 15'h454D: d <= 8'h00; 15'h454E: d <= 8'h00; 15'h454F: d <= 8'h00;
                15'h4550: d <= 8'h00; 15'h4551: d <= 8'h00; 15'h4552: d <= 8'h00; 15'h4553: d <= 8'h00;
                15'h4554: d <= 8'h00; 15'h4555: d <= 8'h00; 15'h4556: d <= 8'h00; 15'h4557: d <= 8'h00;
                15'h4558: d <= 8'h45; 15'h4559: d <= 8'h35; 15'h455A: d <= 8'hAA; 15'h455B: d <= 8'h00;
                15'h455C: d <= 8'h00; 15'h455D: d <= 8'h00; 15'h455E: d <= 8'h00; 15'h455F: d <= 8'h00;
                15'h4560: d <= 8'h00; 15'h4561: d <= 8'h00; 15'h4562: d <= 8'h00; 15'h4563: d <= 8'h00;
                15'h4564: d <= 8'h00; 15'h4565: d <= 8'h00; 15'h4566: d <= 8'h00; 15'h4567: d <= 8'h00;
                15'h4568: d <= 8'h00; 15'h4569: d <= 8'h00; 15'h456A: d <= 8'h00; 15'h456B: d <= 8'h00;
                15'h456C: d <= 8'h00; 15'h456D: d <= 8'h00; 15'h456E: d <= 8'h00; 15'h456F: d <= 8'h00;
                15'h4570: d <= 8'h00; 15'h4571: d <= 8'h00; 15'h4572: d <= 8'h00; 15'h4573: d <= 8'h00;
                15'h4574: d <= 8'h00; 15'h4575: d <= 8'h00; 15'h4576: d <= 8'h00; 15'h4577: d <= 8'h00;
                15'h4578: d <= 8'h00; 15'h4579: d <= 8'h00; 15'h457A: d <= 8'h00; 15'h457B: d <= 8'h00;
                15'h457C: d <= 8'h00; 15'h457D: d <= 8'h00; 15'h457E: d <= 8'h00; 15'h457F: d <= 8'hE0;
                15'h4580: d <= 8'h10; 15'h4581: d <= 8'h15; 15'h4582: d <= 8'h1A; 15'h4583: d <= 8'h1F;
                15'h4584: d <= 8'h20; 15'h4585: d <= 8'h25; 15'h4586: d <= 8'h2A; 15'h4587: d <= 8'h2F;
                15'h4588: d <= 8'h34; 15'h4589: d <= 8'h38; 15'h458A: d <= 8'h3C; 15'h458B: d <= 8'h31;
                15'h458C: d <= 8'h39; 15'h458D: d <= 8'h3D; 15'h458E: d <= 8'h32; 15'h458F: d <= 8'h36;
                15'h4590: d <= 8'h3E; 15'h4591: d <= 8'h33; 15'h4592: d <= 8'h37; 15'h4593: d <= 8'h3B;
                15'h4594: d <= 8'h44; 15'h4595: d <= 8'h48; 15'h4596: d <= 8'h4C; 15'h4597: d <= 8'h41;
                15'h4598: d <= 8'h49; 15'h4599: d <= 8'h4D; 15'h459A: d <= 8'h42; 15'h459B: d <= 8'h46;
                15'h459C: d <= 8'h4E; 15'h459D: d <= 8'h43; 15'h459E: d <= 8'h47; 15'h459F: d <= 8'h4B;
                15'h45A0: d <= 8'h50; 15'h45A1: d <= 8'h55; 15'h45A2: d <= 8'h5A; 15'h45A3: d <= 8'h5F;
                15'h45A4: d <= 8'h60; 15'h45A5: d <= 8'h65; 15'h45A6: d <= 8'h6A; 15'h45A7: d <= 8'h6F;
                15'h45A8: d <= 8'h74; 15'h45A9: d <= 8'h78; 15'h45AA: d <= 8'h7C; 15'h45AB: d <= 8'h71;
                15'h45AC: d <= 8'h79; 15'h45AD: d <= 8'h7D; 15'h45AE: d <= 8'h72; 15'h45AF: d <= 8'h76;
                15'h45B0: d <= 8'h7E; 15'h45B1: d <= 8'h73; 15'h45B2: d <= 8'h77; 15'h45B3: d <= 8'h7B;
                15'h45B4: d <= 8'h84; 15'h45B5: d <= 8'h88; 15'h45B6: d <= 8'h8C; 15'h45B7: d <= 8'h81;
                15'h45B8: d <= 8'h89; 15'h45B9: d <= 8'h8D; 15'h45BA: d <= 8'h82; 15'h45BB: d <= 8'h86;
                15'h45BC: d <= 8'h8E; 15'h45BD: d <= 8'h83; 15'h45BE: d <= 8'h87; 15'h45BF: d <= 8'h8B;
                15'h45C0: d <= 8'h90; 15'h45C1: d <= 8'h95; 15'h45C2: d <= 8'h9A; 15'h45C3: d <= 8'h9F;
                15'h45C4: d <= 8'hA4; 15'h45C5: d <= 8'hA8; 15'h45C6: d <= 8'hAC; 15'h45C7: d <= 8'hA1;
                15'h45C8: d <= 8'hA9; 15'h45C9: d <= 8'hAD; 15'h45CA: d <= 8'hA2; 15'h45CB: d <= 8'hA6;
                15'h45CC: d <= 8'hAE; 15'h45CD: d <= 8'hA3; 15'h45CE: d <= 8'hA7; 15'h45CF: d <= 8'hAB;
                15'h45D0: d <= 8'hB4; 15'h45D1: d <= 8'hB8; 15'h45D2: d <= 8'hBC; 15'h45D3: d <= 8'hB1;
                15'h45D4: d <= 8'hB9; 15'h45D5: d <= 8'hBD; 15'h45D6: d <= 8'hB2; 15'h45D7: d <= 8'hB6;
                15'h45D8: d <= 8'hBE; 15'h45D9: d <= 8'hB3; 15'h45DA: d <= 8'hB7; 15'h45DB: d <= 8'hBB;
                15'h45DC: d <= 8'hC4; 15'h45DD: d <= 8'hC8; 15'h45DE: d <= 8'hCC; 15'h45DF: d <= 8'hC1;
                15'h45E0: d <= 8'hC9; 15'h45E1: d <= 8'hCD; 15'h45E2: d <= 8'hC2; 15'h45E3: d <= 8'hC6;
                15'h45E4: d <= 8'hCE; 15'h45E5: d <= 8'hC3; 15'h45E6: d <= 8'hC7; 15'h45E7: d <= 8'hCB;
                15'h45E8: d <= 8'hC0; 15'h45E9: d <= 8'hC5; 15'h45EA: d <= 8'hCA; 15'h45EB: d <= 8'hCF;
                15'h45EC: d <= 8'hD0; 15'h45ED: d <= 8'hD5; 15'h45EE: d <= 8'hDA; 15'h45EF: d <= 8'hDF;
                15'h45F0: d <= 8'h74; 15'h45F1: d <= 8'h78; 15'h45F2: d <= 8'h7C; 15'h45F3: d <= 8'h71;
                15'h45F4: d <= 8'h79; 15'h45F5: d <= 8'h7D; 15'h45F6: d <= 8'h72; 15'h45F7: d <= 8'h76;
                15'h45F8: d <= 8'h7E; 15'h45F9: d <= 8'h73; 15'h45FA: d <= 8'h77; 15'h45FB: d <= 8'h7B;
                15'h45FC: d <= 8'hA0; 15'h45FD: d <= 8'hA5; 15'h45FE: d <= 8'hAA; 15'h45FF: d <= 8'hAF;
                15'h4600: d <= 8'h00; 15'h4601: d <= 8'h00; 15'h4602: d <= 8'h00; 15'h4603: d <= 8'h00;
                15'h4604: d <= 8'h00; 15'h4605: d <= 8'h00; 15'h4606: d <= 8'h00; 15'h4607: d <= 8'h00;
                15'h4608: d <= 8'h00; 15'h4609: d <= 8'h00; 15'h460A: d <= 8'h00; 15'h460B: d <= 8'h00;
                15'h460C: d <= 8'h00; 15'h460D: d <= 8'h00; 15'h460E: d <= 8'h00; 15'h460F: d <= 8'h00;
                15'h4610: d <= 8'h00; 15'h4611: d <= 8'h00; 15'h4612: d <= 8'h00; 15'h4613: d <= 8'h00;
                15'h4614: d <= 8'h00; 15'h4615: d <= 8'h00; 15'h4616: d <= 8'h00; 15'h4617: d <= 8'h00;
                15'h4618: d <= 8'h00; 15'h4619: d <= 8'h00; 15'h461A: d <= 8'h00; 15'h461B: d <= 8'h00;
                15'h461C: d <= 8'h00; 15'h461D: d <= 8'h00; 15'h461E: d <= 8'h00; 15'h461F: d <= 8'h00;
                15'h4620: d <= 8'h00; 15'h4621: d <= 8'h00; 15'h4622: d <= 8'h00; 15'h4623: d <= 8'h00;
                15'h4624: d <= 8'h00; 15'h4625: d <= 8'h00; 15'h4626: d <= 8'h00; 15'h4627: d <= 8'h00;
                15'h4628: d <= 8'h00; 15'h4629: d <= 8'h00; 15'h462A: d <= 8'h00; 15'h462B: d <= 8'h00;
                15'h462C: d <= 8'h00; 15'h462D: d <= 8'h00; 15'h462E: d <= 8'h00; 15'h462F: d <= 8'hAF;
                15'h4630: d <= 8'h00; 15'h4631: d <= 8'h00; 15'h4632: d <= 8'h00; 15'h4633: d <= 8'h00;
                15'h4634: d <= 8'h00; 15'h4635: d <= 8'h00; 15'h4636: d <= 8'h00; 15'h4637: d <= 8'h00;
                15'h4638: d <= 8'h00; 15'h4639: d <= 8'h00; 15'h463A: d <= 8'h00; 15'h463B: d <= 8'h00;
                15'h463C: d <= 8'h00; 15'h463D: d <= 8'h00; 15'h463E: d <= 8'h00; 15'h463F: d <= 8'h00;
                15'h4640: d <= 8'h00; 15'h4641: d <= 8'h00; 15'h4642: d <= 8'h00; 15'h4643: d <= 8'h00;
                15'h4644: d <= 8'h00; 15'h4645: d <= 8'h00; 15'h4646: d <= 8'h00; 15'h4647: d <= 8'h00;
                15'h4648: d <= 8'h00; 15'h4649: d <= 8'h00; 15'h464A: d <= 8'h00; 15'h464B: d <= 8'h00;
                15'h464C: d <= 8'h00; 15'h464D: d <= 8'h00; 15'h464E: d <= 8'h00; 15'h464F: d <= 8'h00;
                15'h4650: d <= 8'h00; 15'h4651: d <= 8'h00; 15'h4652: d <= 8'h00; 15'h4653: d <= 8'h00;
                15'h4654: d <= 8'h00; 15'h4655: d <= 8'h00; 15'h4656: d <= 8'h00; 15'h4657: d <= 8'h00;
                15'h4658: d <= 8'h45; 15'h4659: d <= 8'h35; 15'h465A: d <= 8'hAA; 15'h465B: d <= 8'h00;
                15'h465C: d <= 8'h00; 15'h465D: d <= 8'h00; 15'h465E: d <= 8'h00; 15'h465F: d <= 8'h00;
                15'h4660: d <= 8'h00; 15'h4661: d <= 8'h00; 15'h4662: d <= 8'h00; 15'h4663: d <= 8'h00;
                15'h4664: d <= 8'h00; 15'h4665: d <= 8'h00; 15'h4666: d <= 8'h00; 15'h4667: d <= 8'h00;
                15'h4668: d <= 8'h00; 15'h4669: d <= 8'h00; 15'h466A: d <= 8'h00; 15'h466B: d <= 8'h00;
                15'h466C: d <= 8'h00; 15'h466D: d <= 8'h00; 15'h466E: d <= 8'h00; 15'h466F: d <= 8'h00;
                15'h4670: d <= 8'h00; 15'h4671: d <= 8'h00; 15'h4672: d <= 8'h00; 15'h4673: d <= 8'h00;
                15'h4674: d <= 8'h00; 15'h4675: d <= 8'h00; 15'h4676: d <= 8'h00; 15'h4677: d <= 8'h00;
                15'h4678: d <= 8'h00; 15'h4679: d <= 8'h00; 15'h467A: d <= 8'h00; 15'h467B: d <= 8'h00;
                15'h467C: d <= 8'h00; 15'h467D: d <= 8'h00; 15'h467E: d <= 8'h00; 15'h467F: d <= 8'hE0;
                15'h4680: d <= 8'h10; 15'h4681: d <= 8'h15; 15'h4682: d <= 8'h1A; 15'h4683: d <= 8'h1F;
                15'h4684: d <= 8'h20; 15'h4685: d <= 8'h25; 15'h4686: d <= 8'h2A; 15'h4687: d <= 8'h2F;
                15'h4688: d <= 8'h34; 15'h4689: d <= 8'h38; 15'h468A: d <= 8'h3C; 15'h468B: d <= 8'h31;
                15'h468C: d <= 8'h39; 15'h468D: d <= 8'h3D; 15'h468E: d <= 8'h32; 15'h468F: d <= 8'h36;
                15'h4690: d <= 8'h3E; 15'h4691: d <= 8'h33; 15'h4692: d <= 8'h37; 15'h4693: d <= 8'h3B;
                15'h4694: d <= 8'h44; 15'h4695: d <= 8'h48; 15'h4696: d <= 8'h4C; 15'h4697: d <= 8'h41;
                15'h4698: d <= 8'h49; 15'h4699: d <= 8'h4D; 15'h469A: d <= 8'h42; 15'h469B: d <= 8'h46;
                15'h469C: d <= 8'h4E; 15'h469D: d <= 8'h43; 15'h469E: d <= 8'h47; 15'h469F: d <= 8'h4B;
                15'h46A0: d <= 8'h50; 15'h46A1: d <= 8'h55; 15'h46A2: d <= 8'h5A; 15'h46A3: d <= 8'h5F;
                15'h46A4: d <= 8'h60; 15'h46A5: d <= 8'h65; 15'h46A6: d <= 8'h6A; 15'h46A7: d <= 8'h6F;
                15'h46A8: d <= 8'h74; 15'h46A9: d <= 8'h78; 15'h46AA: d <= 8'h7C; 15'h46AB: d <= 8'h71;
                15'h46AC: d <= 8'h79; 15'h46AD: d <= 8'h7D; 15'h46AE: d <= 8'h72; 15'h46AF: d <= 8'h76;
                15'h46B0: d <= 8'h7E; 15'h46B1: d <= 8'h73; 15'h46B2: d <= 8'h77; 15'h46B3: d <= 8'h7B;
                15'h46B4: d <= 8'h84; 15'h46B5: d <= 8'h88; 15'h46B6: d <= 8'h8C; 15'h46B7: d <= 8'h81;
                15'h46B8: d <= 8'h89; 15'h46B9: d <= 8'h8D; 15'h46BA: d <= 8'h82; 15'h46BB: d <= 8'h86;
                15'h46BC: d <= 8'h8E; 15'h46BD: d <= 8'h83; 15'h46BE: d <= 8'h87; 15'h46BF: d <= 8'h8B;
                15'h46C0: d <= 8'h90; 15'h46C1: d <= 8'h95; 15'h46C2: d <= 8'h9A; 15'h46C3: d <= 8'h9F;
                15'h46C4: d <= 8'hA4; 15'h46C5: d <= 8'hA8; 15'h46C6: d <= 8'hAC; 15'h46C7: d <= 8'hA1;
                15'h46C8: d <= 8'hA9; 15'h46C9: d <= 8'hAD; 15'h46CA: d <= 8'hA2; 15'h46CB: d <= 8'hA6;
                15'h46CC: d <= 8'hAE; 15'h46CD: d <= 8'hA3; 15'h46CE: d <= 8'hA7; 15'h46CF: d <= 8'hAB;
                15'h46D0: d <= 8'hB4; 15'h46D1: d <= 8'hB8; 15'h46D2: d <= 8'hBC; 15'h46D3: d <= 8'hB1;
                15'h46D4: d <= 8'hB9; 15'h46D5: d <= 8'hBD; 15'h46D6: d <= 8'hB2; 15'h46D7: d <= 8'hB6;
                15'h46D8: d <= 8'hBE; 15'h46D9: d <= 8'hB3; 15'h46DA: d <= 8'hB7; 15'h46DB: d <= 8'hBB;
                15'h46DC: d <= 8'hC4; 15'h46DD: d <= 8'hC8; 15'h46DE: d <= 8'hCC; 15'h46DF: d <= 8'hC1;
                15'h46E0: d <= 8'hC9; 15'h46E1: d <= 8'hCD; 15'h46E2: d <= 8'hC2; 15'h46E3: d <= 8'hC6;
                15'h46E4: d <= 8'hCE; 15'h46E5: d <= 8'hC3; 15'h46E6: d <= 8'hC7; 15'h46E7: d <= 8'hCB;
                15'h46E8: d <= 8'hC0; 15'h46E9: d <= 8'hC5; 15'h46EA: d <= 8'hCA; 15'h46EB: d <= 8'hCF;
                15'h46EC: d <= 8'hD0; 15'h46ED: d <= 8'hD5; 15'h46EE: d <= 8'hDA; 15'h46EF: d <= 8'hDF;
                15'h46F0: d <= 8'h74; 15'h46F1: d <= 8'h78; 15'h46F2: d <= 8'h7C; 15'h46F3: d <= 8'h71;
                15'h46F4: d <= 8'h79; 15'h46F5: d <= 8'h7D; 15'h46F6: d <= 8'h72; 15'h46F7: d <= 8'h76;
                15'h46F8: d <= 8'h7E; 15'h46F9: d <= 8'h73; 15'h46FA: d <= 8'h77; 15'h46FB: d <= 8'h7B;
                15'h46FC: d <= 8'hA0; 15'h46FD: d <= 8'hA5; 15'h46FE: d <= 8'hAA; 15'h46FF: d <= 8'hAF;
                15'h4700: d <= 8'h00; 15'h4701: d <= 8'h00; 15'h4702: d <= 8'h00; 15'h4703: d <= 8'h00;
                15'h4704: d <= 8'h00; 15'h4705: d <= 8'h00; 15'h4706: d <= 8'h00; 15'h4707: d <= 8'h00;
                15'h4708: d <= 8'h00; 15'h4709: d <= 8'h00; 15'h470A: d <= 8'h00; 15'h470B: d <= 8'h00;
                15'h470C: d <= 8'h00; 15'h470D: d <= 8'h00; 15'h470E: d <= 8'h00; 15'h470F: d <= 8'h00;
                15'h4710: d <= 8'h00; 15'h4711: d <= 8'h00; 15'h4712: d <= 8'h00; 15'h4713: d <= 8'h00;
                15'h4714: d <= 8'h00; 15'h4715: d <= 8'h00; 15'h4716: d <= 8'h00; 15'h4717: d <= 8'h00;
                15'h4718: d <= 8'h00; 15'h4719: d <= 8'h00; 15'h471A: d <= 8'h00; 15'h471B: d <= 8'h00;
                15'h471C: d <= 8'h00; 15'h471D: d <= 8'h00; 15'h471E: d <= 8'h00; 15'h471F: d <= 8'h00;
                15'h4720: d <= 8'h00; 15'h4721: d <= 8'h00; 15'h4722: d <= 8'h00; 15'h4723: d <= 8'h00;
                15'h4724: d <= 8'h00; 15'h4725: d <= 8'h00; 15'h4726: d <= 8'h00; 15'h4727: d <= 8'h00;
                15'h4728: d <= 8'h00; 15'h4729: d <= 8'h00; 15'h472A: d <= 8'h00; 15'h472B: d <= 8'h00;
                15'h472C: d <= 8'h00; 15'h472D: d <= 8'h00; 15'h472E: d <= 8'h00; 15'h472F: d <= 8'hAF;
                15'h4730: d <= 8'h00; 15'h4731: d <= 8'h00; 15'h4732: d <= 8'h00; 15'h4733: d <= 8'h00;
                15'h4734: d <= 8'h00; 15'h4735: d <= 8'h00; 15'h4736: d <= 8'h00; 15'h4737: d <= 8'h00;
                15'h4738: d <= 8'h00; 15'h4739: d <= 8'h00; 15'h473A: d <= 8'h00; 15'h473B: d <= 8'h00;
                15'h473C: d <= 8'h00; 15'h473D: d <= 8'h00; 15'h473E: d <= 8'h00; 15'h473F: d <= 8'h00;
                15'h4740: d <= 8'h00; 15'h4741: d <= 8'h00; 15'h4742: d <= 8'h00; 15'h4743: d <= 8'h00;
                15'h4744: d <= 8'h00; 15'h4745: d <= 8'h00; 15'h4746: d <= 8'h00; 15'h4747: d <= 8'h00;
                15'h4748: d <= 8'h00; 15'h4749: d <= 8'h00; 15'h474A: d <= 8'h00; 15'h474B: d <= 8'h00;
                15'h474C: d <= 8'h00; 15'h474D: d <= 8'h00; 15'h474E: d <= 8'h00; 15'h474F: d <= 8'h00;
                15'h4750: d <= 8'h00; 15'h4751: d <= 8'h00; 15'h4752: d <= 8'h00; 15'h4753: d <= 8'h00;
                15'h4754: d <= 8'h00; 15'h4755: d <= 8'h00; 15'h4756: d <= 8'h00; 15'h4757: d <= 8'h00;
                15'h4758: d <= 8'h45; 15'h4759: d <= 8'h35; 15'h475A: d <= 8'hAA; 15'h475B: d <= 8'h00;
                15'h475C: d <= 8'h00; 15'h475D: d <= 8'h00; 15'h475E: d <= 8'h00; 15'h475F: d <= 8'h00;
                15'h4760: d <= 8'h00; 15'h4761: d <= 8'h00; 15'h4762: d <= 8'h00; 15'h4763: d <= 8'h00;
                15'h4764: d <= 8'h00; 15'h4765: d <= 8'h00; 15'h4766: d <= 8'h00; 15'h4767: d <= 8'h00;
                15'h4768: d <= 8'h00; 15'h4769: d <= 8'h00; 15'h476A: d <= 8'h00; 15'h476B: d <= 8'h00;
                15'h476C: d <= 8'h00; 15'h476D: d <= 8'h00; 15'h476E: d <= 8'h00; 15'h476F: d <= 8'h00;
                15'h4770: d <= 8'h00; 15'h4771: d <= 8'h00; 15'h4772: d <= 8'h00; 15'h4773: d <= 8'h00;
                15'h4774: d <= 8'h00; 15'h4775: d <= 8'h00; 15'h4776: d <= 8'h00; 15'h4777: d <= 8'h00;
                15'h4778: d <= 8'h00; 15'h4779: d <= 8'h00; 15'h477A: d <= 8'h00; 15'h477B: d <= 8'h00;
                15'h477C: d <= 8'h00; 15'h477D: d <= 8'h00; 15'h477E: d <= 8'h00; 15'h477F: d <= 8'hE0;
                15'h4780: d <= 8'h10; 15'h4781: d <= 8'h15; 15'h4782: d <= 8'h1A; 15'h4783: d <= 8'h1F;
                15'h4784: d <= 8'h20; 15'h4785: d <= 8'h25; 15'h4786: d <= 8'h2A; 15'h4787: d <= 8'h2F;
                15'h4788: d <= 8'h34; 15'h4789: d <= 8'h38; 15'h478A: d <= 8'h3C; 15'h478B: d <= 8'h31;
                15'h478C: d <= 8'h39; 15'h478D: d <= 8'h3D; 15'h478E: d <= 8'h32; 15'h478F: d <= 8'h36;
                15'h4790: d <= 8'h3E; 15'h4791: d <= 8'h33; 15'h4792: d <= 8'h37; 15'h4793: d <= 8'h3B;
                15'h4794: d <= 8'h44; 15'h4795: d <= 8'h48; 15'h4796: d <= 8'h4C; 15'h4797: d <= 8'h41;
                15'h4798: d <= 8'h49; 15'h4799: d <= 8'h4D; 15'h479A: d <= 8'h42; 15'h479B: d <= 8'h46;
                15'h479C: d <= 8'h4E; 15'h479D: d <= 8'h43; 15'h479E: d <= 8'h47; 15'h479F: d <= 8'h4B;
                15'h47A0: d <= 8'h50; 15'h47A1: d <= 8'h55; 15'h47A2: d <= 8'h5A; 15'h47A3: d <= 8'h5F;
                15'h47A4: d <= 8'h60; 15'h47A5: d <= 8'h65; 15'h47A6: d <= 8'h6A; 15'h47A7: d <= 8'h6F;
                15'h47A8: d <= 8'h74; 15'h47A9: d <= 8'h78; 15'h47AA: d <= 8'h7C; 15'h47AB: d <= 8'h71;
                15'h47AC: d <= 8'h79; 15'h47AD: d <= 8'h7D; 15'h47AE: d <= 8'h72; 15'h47AF: d <= 8'h76;
                15'h47B0: d <= 8'h7E; 15'h47B1: d <= 8'h73; 15'h47B2: d <= 8'h77; 15'h47B3: d <= 8'h7B;
                15'h47B4: d <= 8'h84; 15'h47B5: d <= 8'h88; 15'h47B6: d <= 8'h8C; 15'h47B7: d <= 8'h81;
                15'h47B8: d <= 8'h89; 15'h47B9: d <= 8'h8D; 15'h47BA: d <= 8'h82; 15'h47BB: d <= 8'h86;
                15'h47BC: d <= 8'h8E; 15'h47BD: d <= 8'h83; 15'h47BE: d <= 8'h87; 15'h47BF: d <= 8'h8B;
                15'h47C0: d <= 8'h90; 15'h47C1: d <= 8'h95; 15'h47C2: d <= 8'h9A; 15'h47C3: d <= 8'h9F;
                15'h47C4: d <= 8'hA4; 15'h47C5: d <= 8'hA8; 15'h47C6: d <= 8'hAC; 15'h47C7: d <= 8'hA1;
                15'h47C8: d <= 8'hA9; 15'h47C9: d <= 8'hAD; 15'h47CA: d <= 8'hA2; 15'h47CB: d <= 8'hA6;
                15'h47CC: d <= 8'hAE; 15'h47CD: d <= 8'hA3; 15'h47CE: d <= 8'hA7; 15'h47CF: d <= 8'hAB;
                15'h47D0: d <= 8'hB4; 15'h47D1: d <= 8'hB8; 15'h47D2: d <= 8'hBC; 15'h47D3: d <= 8'hB1;
                15'h47D4: d <= 8'hB9; 15'h47D5: d <= 8'hBD; 15'h47D6: d <= 8'hB2; 15'h47D7: d <= 8'hB6;
                15'h47D8: d <= 8'hBE; 15'h47D9: d <= 8'hB3; 15'h47DA: d <= 8'hB7; 15'h47DB: d <= 8'hBB;
                15'h47DC: d <= 8'hC4; 15'h47DD: d <= 8'hC8; 15'h47DE: d <= 8'hCC; 15'h47DF: d <= 8'hC1;
                15'h47E0: d <= 8'hC9; 15'h47E1: d <= 8'hCD; 15'h47E2: d <= 8'hC2; 15'h47E3: d <= 8'hC6;
                15'h47E4: d <= 8'hCE; 15'h47E5: d <= 8'hC3; 15'h47E6: d <= 8'hC7; 15'h47E7: d <= 8'hCB;
                15'h47E8: d <= 8'hC0; 15'h47E9: d <= 8'hC5; 15'h47EA: d <= 8'hCA; 15'h47EB: d <= 8'hCF;
                15'h47EC: d <= 8'hD0; 15'h47ED: d <= 8'hD5; 15'h47EE: d <= 8'hDA; 15'h47EF: d <= 8'hDF;
                15'h47F0: d <= 8'h74; 15'h47F1: d <= 8'h78; 15'h47F2: d <= 8'h7C; 15'h47F3: d <= 8'h71;
                15'h47F4: d <= 8'h79; 15'h47F5: d <= 8'h7D; 15'h47F6: d <= 8'h72; 15'h47F7: d <= 8'h76;
                15'h47F8: d <= 8'h7E; 15'h47F9: d <= 8'h73; 15'h47FA: d <= 8'h77; 15'h47FB: d <= 8'h7B;
                15'h47FC: d <= 8'hA0; 15'h47FD: d <= 8'hA5; 15'h47FE: d <= 8'hAA; 15'h47FF: d <= 8'hAF;
                15'h4800: d <= 8'h00; 15'h4801: d <= 8'h00; 15'h4802: d <= 8'h00; 15'h4803: d <= 8'h00;
                15'h4804: d <= 8'h00; 15'h4805: d <= 8'h00; 15'h4806: d <= 8'h00; 15'h4807: d <= 8'h00;
                15'h4808: d <= 8'h00; 15'h4809: d <= 8'h00; 15'h480A: d <= 8'h00; 15'h480B: d <= 8'h00;
                15'h480C: d <= 8'h00; 15'h480D: d <= 8'h00; 15'h480E: d <= 8'h00; 15'h480F: d <= 8'h00;
                15'h4810: d <= 8'h00; 15'h4811: d <= 8'h00; 15'h4812: d <= 8'h00; 15'h4813: d <= 8'h00;
                15'h4814: d <= 8'h00; 15'h4815: d <= 8'h00; 15'h4816: d <= 8'h00; 15'h4817: d <= 8'h00;
                15'h4818: d <= 8'h00; 15'h4819: d <= 8'h00; 15'h481A: d <= 8'h00; 15'h481B: d <= 8'h00;
                15'h481C: d <= 8'h00; 15'h481D: d <= 8'h00; 15'h481E: d <= 8'h00; 15'h481F: d <= 8'h00;
                15'h4820: d <= 8'h00; 15'h4821: d <= 8'h00; 15'h4822: d <= 8'h00; 15'h4823: d <= 8'h00;
                15'h4824: d <= 8'h00; 15'h4825: d <= 8'h00; 15'h4826: d <= 8'h00; 15'h4827: d <= 8'h00;
                15'h4828: d <= 8'h00; 15'h4829: d <= 8'h00; 15'h482A: d <= 8'h00; 15'h482B: d <= 8'h00;
                15'h482C: d <= 8'h00; 15'h482D: d <= 8'h00; 15'h482E: d <= 8'h00; 15'h482F: d <= 8'h7B;
                15'h4830: d <= 8'h00; 15'h4831: d <= 8'h00; 15'h4832: d <= 8'h00; 15'h4833: d <= 8'h00;
                15'h4834: d <= 8'h00; 15'h4835: d <= 8'h00; 15'h4836: d <= 8'h00; 15'h4837: d <= 8'h00;
                15'h4838: d <= 8'h00; 15'h4839: d <= 8'h00; 15'h483A: d <= 8'h00; 15'h483B: d <= 8'h00;
                15'h483C: d <= 8'h00; 15'h483D: d <= 8'h00; 15'h483E: d <= 8'h00; 15'h483F: d <= 8'h00;
                15'h4840: d <= 8'h00; 15'h4841: d <= 8'h00; 15'h4842: d <= 8'h00; 15'h4843: d <= 8'h00;
                15'h4844: d <= 8'h00; 15'h4845: d <= 8'h00; 15'h4846: d <= 8'h00; 15'h4847: d <= 8'h00;
                15'h4848: d <= 8'h00; 15'h4849: d <= 8'h00; 15'h484A: d <= 8'h00; 15'h484B: d <= 8'h00;
                15'h484C: d <= 8'h00; 15'h484D: d <= 8'h00; 15'h484E: d <= 8'h00; 15'h484F: d <= 8'h00;
                15'h4850: d <= 8'h00; 15'h4851: d <= 8'h00; 15'h4852: d <= 8'h00; 15'h4853: d <= 8'h00;
                15'h4854: d <= 8'h00; 15'h4855: d <= 8'h00; 15'h4856: d <= 8'h00; 15'h4857: d <= 8'h00;
                15'h4858: d <= 8'h45; 15'h4859: d <= 8'h35; 15'h485A: d <= 8'h32; 15'h485B: d <= 8'h00;
                15'h485C: d <= 8'h00; 15'h485D: d <= 8'h00; 15'h485E: d <= 8'h00; 15'h485F: d <= 8'h00;
                15'h4860: d <= 8'h00; 15'h4861: d <= 8'h00; 15'h4862: d <= 8'h00; 15'h4863: d <= 8'h00;
                15'h4864: d <= 8'h00; 15'h4865: d <= 8'h00; 15'h4866: d <= 8'h00; 15'h4867: d <= 8'h00;
                15'h4868: d <= 8'h00; 15'h4869: d <= 8'h00; 15'h486A: d <= 8'h00; 15'h486B: d <= 8'h00;
                15'h486C: d <= 8'h00; 15'h486D: d <= 8'h00; 15'h486E: d <= 8'h00; 15'h486F: d <= 8'h00;
                15'h4870: d <= 8'h00; 15'h4871: d <= 8'h00; 15'h4872: d <= 8'h00; 15'h4873: d <= 8'h00;
                15'h4874: d <= 8'h00; 15'h4875: d <= 8'h00; 15'h4876: d <= 8'h00; 15'h4877: d <= 8'h00;
                15'h4878: d <= 8'h00; 15'h4879: d <= 8'h00; 15'h487A: d <= 8'h00; 15'h487B: d <= 8'h00;
                15'h487C: d <= 8'h00; 15'h487D: d <= 8'h00; 15'h487E: d <= 8'h00; 15'h487F: d <= 8'hE0;
                15'h4880: d <= 8'h10; 15'h4881: d <= 8'h15; 15'h4882: d <= 8'h1A; 15'h4883: d <= 8'h1F;
                15'h4884: d <= 8'h20; 15'h4885: d <= 8'h25; 15'h4886: d <= 8'h2A; 15'h4887: d <= 8'h2F;
                15'h4888: d <= 8'h34; 15'h4889: d <= 8'h38; 15'h488A: d <= 8'h3C; 15'h488B: d <= 8'h31;
                15'h488C: d <= 8'h39; 15'h488D: d <= 8'h3D; 15'h488E: d <= 8'h32; 15'h488F: d <= 8'h36;
                15'h4890: d <= 8'h3E; 15'h4891: d <= 8'h33; 15'h4892: d <= 8'h37; 15'h4893: d <= 8'h3B;
                15'h4894: d <= 8'h44; 15'h4895: d <= 8'h48; 15'h4896: d <= 8'h4C; 15'h4897: d <= 8'h41;
                15'h4898: d <= 8'h49; 15'h4899: d <= 8'h4D; 15'h489A: d <= 8'h42; 15'h489B: d <= 8'h46;
                15'h489C: d <= 8'h4E; 15'h489D: d <= 8'h43; 15'h489E: d <= 8'h47; 15'h489F: d <= 8'h4B;
                15'h48A0: d <= 8'h50; 15'h48A1: d <= 8'h55; 15'h48A2: d <= 8'h5A; 15'h48A3: d <= 8'h5F;
                15'h48A4: d <= 8'h60; 15'h48A5: d <= 8'h65; 15'h48A6: d <= 8'h6A; 15'h48A7: d <= 8'h6F;
                15'h48A8: d <= 8'h74; 15'h48A9: d <= 8'h78; 15'h48AA: d <= 8'h7C; 15'h48AB: d <= 8'h71;
                15'h48AC: d <= 8'h79; 15'h48AD: d <= 8'h7D; 15'h48AE: d <= 8'h72; 15'h48AF: d <= 8'h76;
                15'h48B0: d <= 8'h7E; 15'h48B1: d <= 8'h73; 15'h48B2: d <= 8'h77; 15'h48B3: d <= 8'h7B;
                15'h48B4: d <= 8'h84; 15'h48B5: d <= 8'h88; 15'h48B6: d <= 8'h8C; 15'h48B7: d <= 8'h81;
                15'h48B8: d <= 8'h89; 15'h48B9: d <= 8'h8D; 15'h48BA: d <= 8'h82; 15'h48BB: d <= 8'h86;
                15'h48BC: d <= 8'h8E; 15'h48BD: d <= 8'h83; 15'h48BE: d <= 8'h87; 15'h48BF: d <= 8'h8B;
                15'h48C0: d <= 8'h90; 15'h48C1: d <= 8'h95; 15'h48C2: d <= 8'h9A; 15'h48C3: d <= 8'h9F;
                15'h48C4: d <= 8'hA4; 15'h48C5: d <= 8'hA8; 15'h48C6: d <= 8'hAC; 15'h48C7: d <= 8'hA1;
                15'h48C8: d <= 8'hA9; 15'h48C9: d <= 8'hAD; 15'h48CA: d <= 8'hA2; 15'h48CB: d <= 8'hA6;
                15'h48CC: d <= 8'hAE; 15'h48CD: d <= 8'hA3; 15'h48CE: d <= 8'hA7; 15'h48CF: d <= 8'hAB;
                15'h48D0: d <= 8'hB4; 15'h48D1: d <= 8'hB8; 15'h48D2: d <= 8'hBC; 15'h48D3: d <= 8'hB1;
                15'h48D4: d <= 8'hB9; 15'h48D5: d <= 8'hBD; 15'h48D6: d <= 8'hB2; 15'h48D7: d <= 8'hB6;
                15'h48D8: d <= 8'hBE; 15'h48D9: d <= 8'hB3; 15'h48DA: d <= 8'hB7; 15'h48DB: d <= 8'hBB;
                15'h48DC: d <= 8'hC4; 15'h48DD: d <= 8'hC8; 15'h48DE: d <= 8'hCC; 15'h48DF: d <= 8'hC1;
                15'h48E0: d <= 8'hC9; 15'h48E1: d <= 8'hCD; 15'h48E2: d <= 8'hC2; 15'h48E3: d <= 8'hC6;
                15'h48E4: d <= 8'hCE; 15'h48E5: d <= 8'hC3; 15'h48E6: d <= 8'hC7; 15'h48E7: d <= 8'hCB;
                15'h48E8: d <= 8'hC0; 15'h48E9: d <= 8'hC5; 15'h48EA: d <= 8'hCA; 15'h48EB: d <= 8'hCF;
                15'h48EC: d <= 8'hD0; 15'h48ED: d <= 8'hD5; 15'h48EE: d <= 8'hDA; 15'h48EF: d <= 8'hDF;
                15'h48F0: d <= 8'h74; 15'h48F1: d <= 8'h78; 15'h48F2: d <= 8'h7C; 15'h48F3: d <= 8'h71;
                15'h48F4: d <= 8'h79; 15'h48F5: d <= 8'h7D; 15'h48F6: d <= 8'h72; 15'h48F7: d <= 8'h76;
                15'h48F8: d <= 8'h7E; 15'h48F9: d <= 8'h73; 15'h48FA: d <= 8'h77; 15'h48FB: d <= 8'h7B;
                15'h48FC: d <= 8'hA0; 15'h48FD: d <= 8'hA5; 15'h48FE: d <= 8'hAA; 15'h48FF: d <= 8'hAF;
                15'h4900: d <= 8'h00; 15'h4901: d <= 8'h00; 15'h4902: d <= 8'h00; 15'h4903: d <= 8'h00;
                15'h4904: d <= 8'h00; 15'h4905: d <= 8'h00; 15'h4906: d <= 8'h00; 15'h4907: d <= 8'h00;
                15'h4908: d <= 8'h00; 15'h4909: d <= 8'h00; 15'h490A: d <= 8'h00; 15'h490B: d <= 8'h00;
                15'h490C: d <= 8'h00; 15'h490D: d <= 8'h00; 15'h490E: d <= 8'h00; 15'h490F: d <= 8'h00;
                15'h4910: d <= 8'h00; 15'h4911: d <= 8'h00; 15'h4912: d <= 8'h00; 15'h4913: d <= 8'h00;
                15'h4914: d <= 8'h00; 15'h4915: d <= 8'h00; 15'h4916: d <= 8'h00; 15'h4917: d <= 8'h00;
                15'h4918: d <= 8'h00; 15'h4919: d <= 8'h00; 15'h491A: d <= 8'h00; 15'h491B: d <= 8'h00;
                15'h491C: d <= 8'h00; 15'h491D: d <= 8'h00; 15'h491E: d <= 8'h00; 15'h491F: d <= 8'h00;
                15'h4920: d <= 8'h00; 15'h4921: d <= 8'h00; 15'h4922: d <= 8'h00; 15'h4923: d <= 8'h00;
                15'h4924: d <= 8'h00; 15'h4925: d <= 8'h00; 15'h4926: d <= 8'h00; 15'h4927: d <= 8'h00;
                15'h4928: d <= 8'h00; 15'h4929: d <= 8'h00; 15'h492A: d <= 8'h00; 15'h492B: d <= 8'h00;
                15'h492C: d <= 8'h00; 15'h492D: d <= 8'h00; 15'h492E: d <= 8'h00; 15'h492F: d <= 8'h7B;
                15'h4930: d <= 8'h00; 15'h4931: d <= 8'h00; 15'h4932: d <= 8'h00; 15'h4933: d <= 8'h00;
                15'h4934: d <= 8'h00; 15'h4935: d <= 8'h00; 15'h4936: d <= 8'h00; 15'h4937: d <= 8'h00;
                15'h4938: d <= 8'h00; 15'h4939: d <= 8'h00; 15'h493A: d <= 8'h00; 15'h493B: d <= 8'h00;
                15'h493C: d <= 8'h00; 15'h493D: d <= 8'h00; 15'h493E: d <= 8'h00; 15'h493F: d <= 8'h00;
                15'h4940: d <= 8'h00; 15'h4941: d <= 8'h00; 15'h4942: d <= 8'h00; 15'h4943: d <= 8'h00;
                15'h4944: d <= 8'h00; 15'h4945: d <= 8'h00; 15'h4946: d <= 8'h00; 15'h4947: d <= 8'h00;
                15'h4948: d <= 8'h00; 15'h4949: d <= 8'h00; 15'h494A: d <= 8'h00; 15'h494B: d <= 8'h00;
                15'h494C: d <= 8'h00; 15'h494D: d <= 8'h00; 15'h494E: d <= 8'h00; 15'h494F: d <= 8'h00;
                15'h4950: d <= 8'h00; 15'h4951: d <= 8'h00; 15'h4952: d <= 8'h00; 15'h4953: d <= 8'h00;
                15'h4954: d <= 8'h00; 15'h4955: d <= 8'h00; 15'h4956: d <= 8'h00; 15'h4957: d <= 8'h00;
                15'h4958: d <= 8'h45; 15'h4959: d <= 8'h35; 15'h495A: d <= 8'h32; 15'h495B: d <= 8'h00;
                15'h495C: d <= 8'h00; 15'h495D: d <= 8'h00; 15'h495E: d <= 8'h00; 15'h495F: d <= 8'h00;
                15'h4960: d <= 8'h00; 15'h4961: d <= 8'h00; 15'h4962: d <= 8'h00; 15'h4963: d <= 8'h00;
                15'h4964: d <= 8'h00; 15'h4965: d <= 8'h00; 15'h4966: d <= 8'h00; 15'h4967: d <= 8'h00;
                15'h4968: d <= 8'h00; 15'h4969: d <= 8'h00; 15'h496A: d <= 8'h00; 15'h496B: d <= 8'h00;
                15'h496C: d <= 8'h00; 15'h496D: d <= 8'h00; 15'h496E: d <= 8'h00; 15'h496F: d <= 8'h00;
                15'h4970: d <= 8'h00; 15'h4971: d <= 8'h00; 15'h4972: d <= 8'h00; 15'h4973: d <= 8'h00;
                15'h4974: d <= 8'h00; 15'h4975: d <= 8'h00; 15'h4976: d <= 8'h00; 15'h4977: d <= 8'h00;
                15'h4978: d <= 8'h00; 15'h4979: d <= 8'h00; 15'h497A: d <= 8'h00; 15'h497B: d <= 8'h00;
                15'h497C: d <= 8'h00; 15'h497D: d <= 8'h00; 15'h497E: d <= 8'h00; 15'h497F: d <= 8'hE0;
                15'h4980: d <= 8'h10; 15'h4981: d <= 8'h15; 15'h4982: d <= 8'h1A; 15'h4983: d <= 8'h1F;
                15'h4984: d <= 8'h20; 15'h4985: d <= 8'h25; 15'h4986: d <= 8'h2A; 15'h4987: d <= 8'h2F;
                15'h4988: d <= 8'h34; 15'h4989: d <= 8'h38; 15'h498A: d <= 8'h3C; 15'h498B: d <= 8'h31;
                15'h498C: d <= 8'h39; 15'h498D: d <= 8'h3D; 15'h498E: d <= 8'h32; 15'h498F: d <= 8'h36;
                15'h4990: d <= 8'h3E; 15'h4991: d <= 8'h33; 15'h4992: d <= 8'h37; 15'h4993: d <= 8'h3B;
                15'h4994: d <= 8'h44; 15'h4995: d <= 8'h48; 15'h4996: d <= 8'h4C; 15'h4997: d <= 8'h41;
                15'h4998: d <= 8'h49; 15'h4999: d <= 8'h4D; 15'h499A: d <= 8'h42; 15'h499B: d <= 8'h46;
                15'h499C: d <= 8'h4E; 15'h499D: d <= 8'h43; 15'h499E: d <= 8'h47; 15'h499F: d <= 8'h4B;
                15'h49A0: d <= 8'h50; 15'h49A1: d <= 8'h55; 15'h49A2: d <= 8'h5A; 15'h49A3: d <= 8'h5F;
                15'h49A4: d <= 8'h60; 15'h49A5: d <= 8'h65; 15'h49A6: d <= 8'h6A; 15'h49A7: d <= 8'h6F;
                15'h49A8: d <= 8'h74; 15'h49A9: d <= 8'h78; 15'h49AA: d <= 8'h7C; 15'h49AB: d <= 8'h71;
                15'h49AC: d <= 8'h79; 15'h49AD: d <= 8'h7D; 15'h49AE: d <= 8'h72; 15'h49AF: d <= 8'h76;
                15'h49B0: d <= 8'h7E; 15'h49B1: d <= 8'h73; 15'h49B2: d <= 8'h77; 15'h49B3: d <= 8'h7B;
                15'h49B4: d <= 8'h84; 15'h49B5: d <= 8'h88; 15'h49B6: d <= 8'h8C; 15'h49B7: d <= 8'h81;
                15'h49B8: d <= 8'h89; 15'h49B9: d <= 8'h8D; 15'h49BA: d <= 8'h82; 15'h49BB: d <= 8'h86;
                15'h49BC: d <= 8'h8E; 15'h49BD: d <= 8'h83; 15'h49BE: d <= 8'h87; 15'h49BF: d <= 8'h8B;
                15'h49C0: d <= 8'h90; 15'h49C1: d <= 8'h95; 15'h49C2: d <= 8'h9A; 15'h49C3: d <= 8'h9F;
                15'h49C4: d <= 8'hA4; 15'h49C5: d <= 8'hA8; 15'h49C6: d <= 8'hAC; 15'h49C7: d <= 8'hA1;
                15'h49C8: d <= 8'hA9; 15'h49C9: d <= 8'hAD; 15'h49CA: d <= 8'hA2; 15'h49CB: d <= 8'hA6;
                15'h49CC: d <= 8'hAE; 15'h49CD: d <= 8'hA3; 15'h49CE: d <= 8'hA7; 15'h49CF: d <= 8'hAB;
                15'h49D0: d <= 8'hB4; 15'h49D1: d <= 8'hB8; 15'h49D2: d <= 8'hBC; 15'h49D3: d <= 8'hB1;
                15'h49D4: d <= 8'hB9; 15'h49D5: d <= 8'hBD; 15'h49D6: d <= 8'hB2; 15'h49D7: d <= 8'hB6;
                15'h49D8: d <= 8'hBE; 15'h49D9: d <= 8'hB3; 15'h49DA: d <= 8'hB7; 15'h49DB: d <= 8'hBB;
                15'h49DC: d <= 8'hC4; 15'h49DD: d <= 8'hC8; 15'h49DE: d <= 8'hCC; 15'h49DF: d <= 8'hC1;
                15'h49E0: d <= 8'hC9; 15'h49E1: d <= 8'hCD; 15'h49E2: d <= 8'hC2; 15'h49E3: d <= 8'hC6;
                15'h49E4: d <= 8'hCE; 15'h49E5: d <= 8'hC3; 15'h49E6: d <= 8'hC7; 15'h49E7: d <= 8'hCB;
                15'h49E8: d <= 8'hC0; 15'h49E9: d <= 8'hC5; 15'h49EA: d <= 8'hCA; 15'h49EB: d <= 8'hCF;
                15'h49EC: d <= 8'hD0; 15'h49ED: d <= 8'hD5; 15'h49EE: d <= 8'hDA; 15'h49EF: d <= 8'hDF;
                15'h49F0: d <= 8'h74; 15'h49F1: d <= 8'h78; 15'h49F2: d <= 8'h7C; 15'h49F3: d <= 8'h71;
                15'h49F4: d <= 8'h79; 15'h49F5: d <= 8'h7D; 15'h49F6: d <= 8'h72; 15'h49F7: d <= 8'h76;
                15'h49F8: d <= 8'h7E; 15'h49F9: d <= 8'h73; 15'h49FA: d <= 8'h77; 15'h49FB: d <= 8'h7B;
                15'h49FC: d <= 8'hA0; 15'h49FD: d <= 8'hA5; 15'h49FE: d <= 8'hAA; 15'h49FF: d <= 8'hAF;
                15'h4A00: d <= 8'h00; 15'h4A01: d <= 8'h00; 15'h4A02: d <= 8'h00; 15'h4A03: d <= 8'h00;
                15'h4A04: d <= 8'h00; 15'h4A05: d <= 8'h00; 15'h4A06: d <= 8'h00; 15'h4A07: d <= 8'h00;
                15'h4A08: d <= 8'h00; 15'h4A09: d <= 8'h00; 15'h4A0A: d <= 8'h00; 15'h4A0B: d <= 8'h00;
                15'h4A0C: d <= 8'h00; 15'h4A0D: d <= 8'h00; 15'h4A0E: d <= 8'h00; 15'h4A0F: d <= 8'h00;
                15'h4A10: d <= 8'h00; 15'h4A11: d <= 8'h00; 15'h4A12: d <= 8'h00; 15'h4A13: d <= 8'h00;
                15'h4A14: d <= 8'h00; 15'h4A15: d <= 8'h00; 15'h4A16: d <= 8'h00; 15'h4A17: d <= 8'h00;
                15'h4A18: d <= 8'h00; 15'h4A19: d <= 8'h00; 15'h4A1A: d <= 8'h00; 15'h4A1B: d <= 8'h00;
                15'h4A1C: d <= 8'h00; 15'h4A1D: d <= 8'h00; 15'h4A1E: d <= 8'h00; 15'h4A1F: d <= 8'h00;
                15'h4A20: d <= 8'h00; 15'h4A21: d <= 8'h00; 15'h4A22: d <= 8'h00; 15'h4A23: d <= 8'h00;
                15'h4A24: d <= 8'h00; 15'h4A25: d <= 8'h00; 15'h4A26: d <= 8'h00; 15'h4A27: d <= 8'h00;
                15'h4A28: d <= 8'h00; 15'h4A29: d <= 8'h00; 15'h4A2A: d <= 8'h00; 15'h4A2B: d <= 8'h00;
                15'h4A2C: d <= 8'h00; 15'h4A2D: d <= 8'h00; 15'h4A2E: d <= 8'h00; 15'h4A2F: d <= 8'h7B;
                15'h4A30: d <= 8'h00; 15'h4A31: d <= 8'h00; 15'h4A32: d <= 8'h00; 15'h4A33: d <= 8'h00;
                15'h4A34: d <= 8'h00; 15'h4A35: d <= 8'h00; 15'h4A36: d <= 8'h00; 15'h4A37: d <= 8'h00;
                15'h4A38: d <= 8'h00; 15'h4A39: d <= 8'h00; 15'h4A3A: d <= 8'h00; 15'h4A3B: d <= 8'h00;
                15'h4A3C: d <= 8'h00; 15'h4A3D: d <= 8'h00; 15'h4A3E: d <= 8'h00; 15'h4A3F: d <= 8'h00;
                15'h4A40: d <= 8'h00; 15'h4A41: d <= 8'h00; 15'h4A42: d <= 8'h00; 15'h4A43: d <= 8'h00;
                15'h4A44: d <= 8'h00; 15'h4A45: d <= 8'h00; 15'h4A46: d <= 8'h00; 15'h4A47: d <= 8'h00;
                15'h4A48: d <= 8'h00; 15'h4A49: d <= 8'h00; 15'h4A4A: d <= 8'h00; 15'h4A4B: d <= 8'h00;
                15'h4A4C: d <= 8'h00; 15'h4A4D: d <= 8'h00; 15'h4A4E: d <= 8'h00; 15'h4A4F: d <= 8'h00;
                15'h4A50: d <= 8'h00; 15'h4A51: d <= 8'h00; 15'h4A52: d <= 8'h00; 15'h4A53: d <= 8'h00;
                15'h4A54: d <= 8'h00; 15'h4A55: d <= 8'h00; 15'h4A56: d <= 8'h00; 15'h4A57: d <= 8'h00;
                15'h4A58: d <= 8'h45; 15'h4A59: d <= 8'h35; 15'h4A5A: d <= 8'h32; 15'h4A5B: d <= 8'h00;
                15'h4A5C: d <= 8'h00; 15'h4A5D: d <= 8'h00; 15'h4A5E: d <= 8'h00; 15'h4A5F: d <= 8'h00;
                15'h4A60: d <= 8'h00; 15'h4A61: d <= 8'h00; 15'h4A62: d <= 8'h00; 15'h4A63: d <= 8'h00;
                15'h4A64: d <= 8'h00; 15'h4A65: d <= 8'h00; 15'h4A66: d <= 8'h00; 15'h4A67: d <= 8'h00;
                15'h4A68: d <= 8'h00; 15'h4A69: d <= 8'h00; 15'h4A6A: d <= 8'h00; 15'h4A6B: d <= 8'h00;
                15'h4A6C: d <= 8'h00; 15'h4A6D: d <= 8'h00; 15'h4A6E: d <= 8'h00; 15'h4A6F: d <= 8'h00;
                15'h4A70: d <= 8'h00; 15'h4A71: d <= 8'h00; 15'h4A72: d <= 8'h00; 15'h4A73: d <= 8'h00;
                15'h4A74: d <= 8'h00; 15'h4A75: d <= 8'h00; 15'h4A76: d <= 8'h00; 15'h4A77: d <= 8'h00;
                15'h4A78: d <= 8'h00; 15'h4A79: d <= 8'h00; 15'h4A7A: d <= 8'h00; 15'h4A7B: d <= 8'h00;
                15'h4A7C: d <= 8'h00; 15'h4A7D: d <= 8'h00; 15'h4A7E: d <= 8'h00; 15'h4A7F: d <= 8'hE0;
                15'h4A80: d <= 8'h10; 15'h4A81: d <= 8'h15; 15'h4A82: d <= 8'h1A; 15'h4A83: d <= 8'h1F;
                15'h4A84: d <= 8'h20; 15'h4A85: d <= 8'h25; 15'h4A86: d <= 8'h2A; 15'h4A87: d <= 8'h2F;
                15'h4A88: d <= 8'h34; 15'h4A89: d <= 8'h38; 15'h4A8A: d <= 8'h3C; 15'h4A8B: d <= 8'h31;
                15'h4A8C: d <= 8'h39; 15'h4A8D: d <= 8'h3D; 15'h4A8E: d <= 8'h32; 15'h4A8F: d <= 8'h36;
                15'h4A90: d <= 8'h3E; 15'h4A91: d <= 8'h33; 15'h4A92: d <= 8'h37; 15'h4A93: d <= 8'h3B;
                15'h4A94: d <= 8'h44; 15'h4A95: d <= 8'h48; 15'h4A96: d <= 8'h4C; 15'h4A97: d <= 8'h41;
                15'h4A98: d <= 8'h49; 15'h4A99: d <= 8'h4D; 15'h4A9A: d <= 8'h42; 15'h4A9B: d <= 8'h46;
                15'h4A9C: d <= 8'h4E; 15'h4A9D: d <= 8'h43; 15'h4A9E: d <= 8'h47; 15'h4A9F: d <= 8'h4B;
                15'h4AA0: d <= 8'h50; 15'h4AA1: d <= 8'h55; 15'h4AA2: d <= 8'h5A; 15'h4AA3: d <= 8'h5F;
                15'h4AA4: d <= 8'h60; 15'h4AA5: d <= 8'h65; 15'h4AA6: d <= 8'h6A; 15'h4AA7: d <= 8'h6F;
                15'h4AA8: d <= 8'h74; 15'h4AA9: d <= 8'h78; 15'h4AAA: d <= 8'h7C; 15'h4AAB: d <= 8'h71;
                15'h4AAC: d <= 8'h79; 15'h4AAD: d <= 8'h7D; 15'h4AAE: d <= 8'h72; 15'h4AAF: d <= 8'h76;
                15'h4AB0: d <= 8'h7E; 15'h4AB1: d <= 8'h73; 15'h4AB2: d <= 8'h77; 15'h4AB3: d <= 8'h7B;
                15'h4AB4: d <= 8'h84; 15'h4AB5: d <= 8'h88; 15'h4AB6: d <= 8'h8C; 15'h4AB7: d <= 8'h81;
                15'h4AB8: d <= 8'h89; 15'h4AB9: d <= 8'h8D; 15'h4ABA: d <= 8'h82; 15'h4ABB: d <= 8'h86;
                15'h4ABC: d <= 8'h8E; 15'h4ABD: d <= 8'h83; 15'h4ABE: d <= 8'h87; 15'h4ABF: d <= 8'h8B;
                15'h4AC0: d <= 8'h90; 15'h4AC1: d <= 8'h95; 15'h4AC2: d <= 8'h9A; 15'h4AC3: d <= 8'h9F;
                15'h4AC4: d <= 8'hA4; 15'h4AC5: d <= 8'hA8; 15'h4AC6: d <= 8'hAC; 15'h4AC7: d <= 8'hA1;
                15'h4AC8: d <= 8'hA9; 15'h4AC9: d <= 8'hAD; 15'h4ACA: d <= 8'hA2; 15'h4ACB: d <= 8'hA6;
                15'h4ACC: d <= 8'hAE; 15'h4ACD: d <= 8'hA3; 15'h4ACE: d <= 8'hA7; 15'h4ACF: d <= 8'hAB;
                15'h4AD0: d <= 8'hB4; 15'h4AD1: d <= 8'hB8; 15'h4AD2: d <= 8'hBC; 15'h4AD3: d <= 8'hB1;
                15'h4AD4: d <= 8'hB9; 15'h4AD5: d <= 8'hBD; 15'h4AD6: d <= 8'hB2; 15'h4AD7: d <= 8'hB6;
                15'h4AD8: d <= 8'hBE; 15'h4AD9: d <= 8'hB3; 15'h4ADA: d <= 8'hB7; 15'h4ADB: d <= 8'hBB;
                15'h4ADC: d <= 8'hC4; 15'h4ADD: d <= 8'hC8; 15'h4ADE: d <= 8'hCC; 15'h4ADF: d <= 8'hC1;
                15'h4AE0: d <= 8'hC9; 15'h4AE1: d <= 8'hCD; 15'h4AE2: d <= 8'hC2; 15'h4AE3: d <= 8'hC6;
                15'h4AE4: d <= 8'hCE; 15'h4AE5: d <= 8'hC3; 15'h4AE6: d <= 8'hC7; 15'h4AE7: d <= 8'hCB;
                15'h4AE8: d <= 8'hC0; 15'h4AE9: d <= 8'hC5; 15'h4AEA: d <= 8'hCA; 15'h4AEB: d <= 8'hCF;
                15'h4AEC: d <= 8'hD0; 15'h4AED: d <= 8'hD5; 15'h4AEE: d <= 8'hDA; 15'h4AEF: d <= 8'hDF;
                15'h4AF0: d <= 8'h74; 15'h4AF1: d <= 8'h78; 15'h4AF2: d <= 8'h7C; 15'h4AF3: d <= 8'h71;
                15'h4AF4: d <= 8'h79; 15'h4AF5: d <= 8'h7D; 15'h4AF6: d <= 8'h72; 15'h4AF7: d <= 8'h76;
                15'h4AF8: d <= 8'h7E; 15'h4AF9: d <= 8'h73; 15'h4AFA: d <= 8'h77; 15'h4AFB: d <= 8'h7B;
                15'h4AFC: d <= 8'hA0; 15'h4AFD: d <= 8'hA5; 15'h4AFE: d <= 8'hAA; 15'h4AFF: d <= 8'hAF;
                15'h4B00: d <= 8'h00; 15'h4B01: d <= 8'h00; 15'h4B02: d <= 8'h00; 15'h4B03: d <= 8'h00;
                15'h4B04: d <= 8'h00; 15'h4B05: d <= 8'h00; 15'h4B06: d <= 8'h00; 15'h4B07: d <= 8'h00;
                15'h4B08: d <= 8'h00; 15'h4B09: d <= 8'h00; 15'h4B0A: d <= 8'h00; 15'h4B0B: d <= 8'h00;
                15'h4B0C: d <= 8'h00; 15'h4B0D: d <= 8'h00; 15'h4B0E: d <= 8'h00; 15'h4B0F: d <= 8'h00;
                15'h4B10: d <= 8'h00; 15'h4B11: d <= 8'h00; 15'h4B12: d <= 8'h00; 15'h4B13: d <= 8'h00;
                15'h4B14: d <= 8'h00; 15'h4B15: d <= 8'h00; 15'h4B16: d <= 8'h00; 15'h4B17: d <= 8'h00;
                15'h4B18: d <= 8'h00; 15'h4B19: d <= 8'h00; 15'h4B1A: d <= 8'h00; 15'h4B1B: d <= 8'h00;
                15'h4B1C: d <= 8'h00; 15'h4B1D: d <= 8'h00; 15'h4B1E: d <= 8'h00; 15'h4B1F: d <= 8'h00;
                15'h4B20: d <= 8'h00; 15'h4B21: d <= 8'h00; 15'h4B22: d <= 8'h00; 15'h4B23: d <= 8'h00;
                15'h4B24: d <= 8'h00; 15'h4B25: d <= 8'h00; 15'h4B26: d <= 8'h00; 15'h4B27: d <= 8'h00;
                15'h4B28: d <= 8'h00; 15'h4B29: d <= 8'h00; 15'h4B2A: d <= 8'h00; 15'h4B2B: d <= 8'h00;
                15'h4B2C: d <= 8'h00; 15'h4B2D: d <= 8'h00; 15'h4B2E: d <= 8'h00; 15'h4B2F: d <= 8'h7B;
                15'h4B30: d <= 8'h00; 15'h4B31: d <= 8'h00; 15'h4B32: d <= 8'h00; 15'h4B33: d <= 8'h00;
                15'h4B34: d <= 8'h00; 15'h4B35: d <= 8'h00; 15'h4B36: d <= 8'h00; 15'h4B37: d <= 8'h00;
                15'h4B38: d <= 8'h00; 15'h4B39: d <= 8'h00; 15'h4B3A: d <= 8'h00; 15'h4B3B: d <= 8'h00;
                15'h4B3C: d <= 8'h00; 15'h4B3D: d <= 8'h00; 15'h4B3E: d <= 8'h00; 15'h4B3F: d <= 8'h00;
                15'h4B40: d <= 8'h00; 15'h4B41: d <= 8'h00; 15'h4B42: d <= 8'h00; 15'h4B43: d <= 8'h00;
                15'h4B44: d <= 8'h00; 15'h4B45: d <= 8'h00; 15'h4B46: d <= 8'h00; 15'h4B47: d <= 8'h00;
                15'h4B48: d <= 8'h00; 15'h4B49: d <= 8'h00; 15'h4B4A: d <= 8'h00; 15'h4B4B: d <= 8'h00;
                15'h4B4C: d <= 8'h00; 15'h4B4D: d <= 8'h00; 15'h4B4E: d <= 8'h00; 15'h4B4F: d <= 8'h00;
                15'h4B50: d <= 8'h00; 15'h4B51: d <= 8'h00; 15'h4B52: d <= 8'h00; 15'h4B53: d <= 8'h00;
                15'h4B54: d <= 8'h00; 15'h4B55: d <= 8'h00; 15'h4B56: d <= 8'h00; 15'h4B57: d <= 8'h00;
                15'h4B58: d <= 8'h45; 15'h4B59: d <= 8'h35; 15'h4B5A: d <= 8'h32; 15'h4B5B: d <= 8'h00;
                15'h4B5C: d <= 8'h00; 15'h4B5D: d <= 8'h00; 15'h4B5E: d <= 8'h00; 15'h4B5F: d <= 8'h00;
                15'h4B60: d <= 8'h00; 15'h4B61: d <= 8'h00; 15'h4B62: d <= 8'h00; 15'h4B63: d <= 8'h00;
                15'h4B64: d <= 8'h00; 15'h4B65: d <= 8'h00; 15'h4B66: d <= 8'h00; 15'h4B67: d <= 8'h00;
                15'h4B68: d <= 8'h00; 15'h4B69: d <= 8'h00; 15'h4B6A: d <= 8'h00; 15'h4B6B: d <= 8'h00;
                15'h4B6C: d <= 8'h00; 15'h4B6D: d <= 8'h00; 15'h4B6E: d <= 8'h00; 15'h4B6F: d <= 8'h00;
                15'h4B70: d <= 8'h00; 15'h4B71: d <= 8'h00; 15'h4B72: d <= 8'h00; 15'h4B73: d <= 8'h00;
                15'h4B74: d <= 8'h00; 15'h4B75: d <= 8'h00; 15'h4B76: d <= 8'h00; 15'h4B77: d <= 8'h00;
                15'h4B78: d <= 8'h00; 15'h4B79: d <= 8'h00; 15'h4B7A: d <= 8'h00; 15'h4B7B: d <= 8'h00;
                15'h4B7C: d <= 8'h00; 15'h4B7D: d <= 8'h00; 15'h4B7E: d <= 8'h00; 15'h4B7F: d <= 8'hE0;
                15'h4B80: d <= 8'h10; 15'h4B81: d <= 8'h15; 15'h4B82: d <= 8'h1A; 15'h4B83: d <= 8'h1F;
                15'h4B84: d <= 8'h20; 15'h4B85: d <= 8'h25; 15'h4B86: d <= 8'h2A; 15'h4B87: d <= 8'h2F;
                15'h4B88: d <= 8'h34; 15'h4B89: d <= 8'h38; 15'h4B8A: d <= 8'h3C; 15'h4B8B: d <= 8'h31;
                15'h4B8C: d <= 8'h39; 15'h4B8D: d <= 8'h3D; 15'h4B8E: d <= 8'h32; 15'h4B8F: d <= 8'h36;
                15'h4B90: d <= 8'h3E; 15'h4B91: d <= 8'h33; 15'h4B92: d <= 8'h37; 15'h4B93: d <= 8'h3B;
                15'h4B94: d <= 8'h44; 15'h4B95: d <= 8'h48; 15'h4B96: d <= 8'h4C; 15'h4B97: d <= 8'h41;
                15'h4B98: d <= 8'h49; 15'h4B99: d <= 8'h4D; 15'h4B9A: d <= 8'h42; 15'h4B9B: d <= 8'h46;
                15'h4B9C: d <= 8'h4E; 15'h4B9D: d <= 8'h43; 15'h4B9E: d <= 8'h47; 15'h4B9F: d <= 8'h4B;
                15'h4BA0: d <= 8'h50; 15'h4BA1: d <= 8'h55; 15'h4BA2: d <= 8'h5A; 15'h4BA3: d <= 8'h5F;
                15'h4BA4: d <= 8'h60; 15'h4BA5: d <= 8'h65; 15'h4BA6: d <= 8'h6A; 15'h4BA7: d <= 8'h6F;
                15'h4BA8: d <= 8'h74; 15'h4BA9: d <= 8'h78; 15'h4BAA: d <= 8'h7C; 15'h4BAB: d <= 8'h71;
                15'h4BAC: d <= 8'h79; 15'h4BAD: d <= 8'h7D; 15'h4BAE: d <= 8'h72; 15'h4BAF: d <= 8'h76;
                15'h4BB0: d <= 8'h7E; 15'h4BB1: d <= 8'h73; 15'h4BB2: d <= 8'h77; 15'h4BB3: d <= 8'h7B;
                15'h4BB4: d <= 8'h84; 15'h4BB5: d <= 8'h88; 15'h4BB6: d <= 8'h8C; 15'h4BB7: d <= 8'h81;
                15'h4BB8: d <= 8'h89; 15'h4BB9: d <= 8'h8D; 15'h4BBA: d <= 8'h82; 15'h4BBB: d <= 8'h86;
                15'h4BBC: d <= 8'h8E; 15'h4BBD: d <= 8'h83; 15'h4BBE: d <= 8'h87; 15'h4BBF: d <= 8'h8B;
                15'h4BC0: d <= 8'h90; 15'h4BC1: d <= 8'h95; 15'h4BC2: d <= 8'h9A; 15'h4BC3: d <= 8'h9F;
                15'h4BC4: d <= 8'hA4; 15'h4BC5: d <= 8'hA8; 15'h4BC6: d <= 8'hAC; 15'h4BC7: d <= 8'hA1;
                15'h4BC8: d <= 8'hA9; 15'h4BC9: d <= 8'hAD; 15'h4BCA: d <= 8'hA2; 15'h4BCB: d <= 8'hA6;
                15'h4BCC: d <= 8'hAE; 15'h4BCD: d <= 8'hA3; 15'h4BCE: d <= 8'hA7; 15'h4BCF: d <= 8'hAB;
                15'h4BD0: d <= 8'hB4; 15'h4BD1: d <= 8'hB8; 15'h4BD2: d <= 8'hBC; 15'h4BD3: d <= 8'hB1;
                15'h4BD4: d <= 8'hB9; 15'h4BD5: d <= 8'hBD; 15'h4BD6: d <= 8'hB2; 15'h4BD7: d <= 8'hB6;
                15'h4BD8: d <= 8'hBE; 15'h4BD9: d <= 8'hB3; 15'h4BDA: d <= 8'hB7; 15'h4BDB: d <= 8'hBB;
                15'h4BDC: d <= 8'hC4; 15'h4BDD: d <= 8'hC8; 15'h4BDE: d <= 8'hCC; 15'h4BDF: d <= 8'hC1;
                15'h4BE0: d <= 8'hC9; 15'h4BE1: d <= 8'hCD; 15'h4BE2: d <= 8'hC2; 15'h4BE3: d <= 8'hC6;
                15'h4BE4: d <= 8'hCE; 15'h4BE5: d <= 8'hC3; 15'h4BE6: d <= 8'hC7; 15'h4BE7: d <= 8'hCB;
                15'h4BE8: d <= 8'hC0; 15'h4BE9: d <= 8'hC5; 15'h4BEA: d <= 8'hCA; 15'h4BEB: d <= 8'hCF;
                15'h4BEC: d <= 8'hD0; 15'h4BED: d <= 8'hD5; 15'h4BEE: d <= 8'hDA; 15'h4BEF: d <= 8'hDF;
                15'h4BF0: d <= 8'h74; 15'h4BF1: d <= 8'h78; 15'h4BF2: d <= 8'h7C; 15'h4BF3: d <= 8'h71;
                15'h4BF4: d <= 8'h79; 15'h4BF5: d <= 8'h7D; 15'h4BF6: d <= 8'h72; 15'h4BF7: d <= 8'h76;
                15'h4BF8: d <= 8'h7E; 15'h4BF9: d <= 8'h73; 15'h4BFA: d <= 8'h77; 15'h4BFB: d <= 8'h7B;
                15'h4BFC: d <= 8'hA0; 15'h4BFD: d <= 8'hA5; 15'h4BFE: d <= 8'hAA; 15'h4BFF: d <= 8'hAF;
                15'h4C00: d <= 8'h00; 15'h4C01: d <= 8'h00; 15'h4C02: d <= 8'h00; 15'h4C03: d <= 8'h00;
                15'h4C04: d <= 8'h00; 15'h4C05: d <= 8'h00; 15'h4C06: d <= 8'h00; 15'h4C07: d <= 8'h00;
                15'h4C08: d <= 8'h00; 15'h4C09: d <= 8'h00; 15'h4C0A: d <= 8'h00; 15'h4C0B: d <= 8'h00;
                15'h4C0C: d <= 8'h00; 15'h4C0D: d <= 8'h00; 15'h4C0E: d <= 8'h00; 15'h4C0F: d <= 8'h00;
                15'h4C10: d <= 8'h00; 15'h4C11: d <= 8'h00; 15'h4C12: d <= 8'h00; 15'h4C13: d <= 8'h00;
                15'h4C14: d <= 8'h00; 15'h4C15: d <= 8'h00; 15'h4C16: d <= 8'h00; 15'h4C17: d <= 8'h00;
                15'h4C18: d <= 8'h00; 15'h4C19: d <= 8'h00; 15'h4C1A: d <= 8'h00; 15'h4C1B: d <= 8'h00;
                15'h4C1C: d <= 8'h00; 15'h4C1D: d <= 8'h00; 15'h4C1E: d <= 8'h00; 15'h4C1F: d <= 8'h00;
                15'h4C20: d <= 8'h00; 15'h4C21: d <= 8'h00; 15'h4C22: d <= 8'h00; 15'h4C23: d <= 8'h00;
                15'h4C24: d <= 8'h00; 15'h4C25: d <= 8'h00; 15'h4C26: d <= 8'h00; 15'h4C27: d <= 8'h00;
                15'h4C28: d <= 8'h00; 15'h4C29: d <= 8'h00; 15'h4C2A: d <= 8'h00; 15'h4C2B: d <= 8'h00;
                15'h4C2C: d <= 8'h00; 15'h4C2D: d <= 8'h00; 15'h4C2E: d <= 8'h00; 15'h4C2F: d <= 8'h7B;
                15'h4C30: d <= 8'h00; 15'h4C31: d <= 8'h00; 15'h4C32: d <= 8'h00; 15'h4C33: d <= 8'h00;
                15'h4C34: d <= 8'h00; 15'h4C35: d <= 8'h00; 15'h4C36: d <= 8'h00; 15'h4C37: d <= 8'h00;
                15'h4C38: d <= 8'h00; 15'h4C39: d <= 8'h00; 15'h4C3A: d <= 8'h00; 15'h4C3B: d <= 8'h00;
                15'h4C3C: d <= 8'h00; 15'h4C3D: d <= 8'h00; 15'h4C3E: d <= 8'h00; 15'h4C3F: d <= 8'h00;
                15'h4C40: d <= 8'h00; 15'h4C41: d <= 8'h00; 15'h4C42: d <= 8'h00; 15'h4C43: d <= 8'h00;
                15'h4C44: d <= 8'h00; 15'h4C45: d <= 8'h00; 15'h4C46: d <= 8'h00; 15'h4C47: d <= 8'h00;
                15'h4C48: d <= 8'h00; 15'h4C49: d <= 8'h00; 15'h4C4A: d <= 8'h00; 15'h4C4B: d <= 8'h00;
                15'h4C4C: d <= 8'h00; 15'h4C4D: d <= 8'h00; 15'h4C4E: d <= 8'h00; 15'h4C4F: d <= 8'h00;
                15'h4C50: d <= 8'h00; 15'h4C51: d <= 8'h00; 15'h4C52: d <= 8'h00; 15'h4C53: d <= 8'h00;
                15'h4C54: d <= 8'h00; 15'h4C55: d <= 8'h00; 15'h4C56: d <= 8'h00; 15'h4C57: d <= 8'h00;
                15'h4C58: d <= 8'h45; 15'h4C59: d <= 8'h35; 15'h4C5A: d <= 8'h32; 15'h4C5B: d <= 8'h00;
                15'h4C5C: d <= 8'h00; 15'h4C5D: d <= 8'h00; 15'h4C5E: d <= 8'h00; 15'h4C5F: d <= 8'h00;
                15'h4C60: d <= 8'h00; 15'h4C61: d <= 8'h00; 15'h4C62: d <= 8'h00; 15'h4C63: d <= 8'h00;
                15'h4C64: d <= 8'h00; 15'h4C65: d <= 8'h00; 15'h4C66: d <= 8'h00; 15'h4C67: d <= 8'h00;
                15'h4C68: d <= 8'h00; 15'h4C69: d <= 8'h00; 15'h4C6A: d <= 8'h00; 15'h4C6B: d <= 8'h00;
                15'h4C6C: d <= 8'h00; 15'h4C6D: d <= 8'h00; 15'h4C6E: d <= 8'h00; 15'h4C6F: d <= 8'h00;
                15'h4C70: d <= 8'h00; 15'h4C71: d <= 8'h00; 15'h4C72: d <= 8'h00; 15'h4C73: d <= 8'h00;
                15'h4C74: d <= 8'h00; 15'h4C75: d <= 8'h00; 15'h4C76: d <= 8'h00; 15'h4C77: d <= 8'h00;
                15'h4C78: d <= 8'h00; 15'h4C79: d <= 8'h00; 15'h4C7A: d <= 8'h00; 15'h4C7B: d <= 8'h00;
                15'h4C7C: d <= 8'h00; 15'h4C7D: d <= 8'h00; 15'h4C7E: d <= 8'h00; 15'h4C7F: d <= 8'hE0;
                15'h4C80: d <= 8'h10; 15'h4C81: d <= 8'h15; 15'h4C82: d <= 8'h1A; 15'h4C83: d <= 8'h1F;
                15'h4C84: d <= 8'h20; 15'h4C85: d <= 8'h25; 15'h4C86: d <= 8'h2A; 15'h4C87: d <= 8'h2F;
                15'h4C88: d <= 8'h34; 15'h4C89: d <= 8'h38; 15'h4C8A: d <= 8'h3C; 15'h4C8B: d <= 8'h31;
                15'h4C8C: d <= 8'h39; 15'h4C8D: d <= 8'h3D; 15'h4C8E: d <= 8'h32; 15'h4C8F: d <= 8'h36;
                15'h4C90: d <= 8'h3E; 15'h4C91: d <= 8'h33; 15'h4C92: d <= 8'h37; 15'h4C93: d <= 8'h3B;
                15'h4C94: d <= 8'h44; 15'h4C95: d <= 8'h48; 15'h4C96: d <= 8'h4C; 15'h4C97: d <= 8'h41;
                15'h4C98: d <= 8'h49; 15'h4C99: d <= 8'h4D; 15'h4C9A: d <= 8'h42; 15'h4C9B: d <= 8'h46;
                15'h4C9C: d <= 8'h4E; 15'h4C9D: d <= 8'h43; 15'h4C9E: d <= 8'h47; 15'h4C9F: d <= 8'h4B;
                15'h4CA0: d <= 8'h50; 15'h4CA1: d <= 8'h55; 15'h4CA2: d <= 8'h5A; 15'h4CA3: d <= 8'h5F;
                15'h4CA4: d <= 8'h60; 15'h4CA5: d <= 8'h65; 15'h4CA6: d <= 8'h6A; 15'h4CA7: d <= 8'h6F;
                15'h4CA8: d <= 8'h74; 15'h4CA9: d <= 8'h78; 15'h4CAA: d <= 8'h7C; 15'h4CAB: d <= 8'h71;
                15'h4CAC: d <= 8'h79; 15'h4CAD: d <= 8'h7D; 15'h4CAE: d <= 8'h72; 15'h4CAF: d <= 8'h76;
                15'h4CB0: d <= 8'h7E; 15'h4CB1: d <= 8'h73; 15'h4CB2: d <= 8'h77; 15'h4CB3: d <= 8'h7B;
                15'h4CB4: d <= 8'h84; 15'h4CB5: d <= 8'h88; 15'h4CB6: d <= 8'h8C; 15'h4CB7: d <= 8'h81;
                15'h4CB8: d <= 8'h89; 15'h4CB9: d <= 8'h8D; 15'h4CBA: d <= 8'h82; 15'h4CBB: d <= 8'h86;
                15'h4CBC: d <= 8'h8E; 15'h4CBD: d <= 8'h83; 15'h4CBE: d <= 8'h87; 15'h4CBF: d <= 8'h8B;
                15'h4CC0: d <= 8'h90; 15'h4CC1: d <= 8'h95; 15'h4CC2: d <= 8'h9A; 15'h4CC3: d <= 8'h9F;
                15'h4CC4: d <= 8'hA4; 15'h4CC5: d <= 8'hA8; 15'h4CC6: d <= 8'hAC; 15'h4CC7: d <= 8'hA1;
                15'h4CC8: d <= 8'hA9; 15'h4CC9: d <= 8'hAD; 15'h4CCA: d <= 8'hA2; 15'h4CCB: d <= 8'hA6;
                15'h4CCC: d <= 8'hAE; 15'h4CCD: d <= 8'hA3; 15'h4CCE: d <= 8'hA7; 15'h4CCF: d <= 8'hAB;
                15'h4CD0: d <= 8'hB4; 15'h4CD1: d <= 8'hB8; 15'h4CD2: d <= 8'hBC; 15'h4CD3: d <= 8'hB1;
                15'h4CD4: d <= 8'hB9; 15'h4CD5: d <= 8'hBD; 15'h4CD6: d <= 8'hB2; 15'h4CD7: d <= 8'hB6;
                15'h4CD8: d <= 8'hBE; 15'h4CD9: d <= 8'hB3; 15'h4CDA: d <= 8'hB7; 15'h4CDB: d <= 8'hBB;
                15'h4CDC: d <= 8'hC4; 15'h4CDD: d <= 8'hC8; 15'h4CDE: d <= 8'hCC; 15'h4CDF: d <= 8'hC1;
                15'h4CE0: d <= 8'hC9; 15'h4CE1: d <= 8'hCD; 15'h4CE2: d <= 8'hC2; 15'h4CE3: d <= 8'hC6;
                15'h4CE4: d <= 8'hCE; 15'h4CE5: d <= 8'hC3; 15'h4CE6: d <= 8'hC7; 15'h4CE7: d <= 8'hCB;
                15'h4CE8: d <= 8'hC0; 15'h4CE9: d <= 8'hC5; 15'h4CEA: d <= 8'hCA; 15'h4CEB: d <= 8'hCF;
                15'h4CEC: d <= 8'hD0; 15'h4CED: d <= 8'hD5; 15'h4CEE: d <= 8'hDA; 15'h4CEF: d <= 8'hDF;
                15'h4CF0: d <= 8'h74; 15'h4CF1: d <= 8'h78; 15'h4CF2: d <= 8'h7C; 15'h4CF3: d <= 8'h71;
                15'h4CF4: d <= 8'h79; 15'h4CF5: d <= 8'h7D; 15'h4CF6: d <= 8'h72; 15'h4CF7: d <= 8'h76;
                15'h4CF8: d <= 8'h7E; 15'h4CF9: d <= 8'h73; 15'h4CFA: d <= 8'h77; 15'h4CFB: d <= 8'h7B;
                15'h4CFC: d <= 8'hA0; 15'h4CFD: d <= 8'hA5; 15'h4CFE: d <= 8'hAA; 15'h4CFF: d <= 8'hAF;
                15'h4D00: d <= 8'h00; 15'h4D01: d <= 8'h00; 15'h4D02: d <= 8'h00; 15'h4D03: d <= 8'h00;
                15'h4D04: d <= 8'h00; 15'h4D05: d <= 8'h00; 15'h4D06: d <= 8'h00; 15'h4D07: d <= 8'h00;
                15'h4D08: d <= 8'h00; 15'h4D09: d <= 8'h00; 15'h4D0A: d <= 8'h00; 15'h4D0B: d <= 8'h00;
                15'h4D0C: d <= 8'h00; 15'h4D0D: d <= 8'h00; 15'h4D0E: d <= 8'h00; 15'h4D0F: d <= 8'h00;
                15'h4D10: d <= 8'h00; 15'h4D11: d <= 8'h00; 15'h4D12: d <= 8'h00; 15'h4D13: d <= 8'h00;
                15'h4D14: d <= 8'h00; 15'h4D15: d <= 8'h00; 15'h4D16: d <= 8'h00; 15'h4D17: d <= 8'h00;
                15'h4D18: d <= 8'h00; 15'h4D19: d <= 8'h00; 15'h4D1A: d <= 8'h00; 15'h4D1B: d <= 8'h00;
                15'h4D1C: d <= 8'h00; 15'h4D1D: d <= 8'h00; 15'h4D1E: d <= 8'h00; 15'h4D1F: d <= 8'h00;
                15'h4D20: d <= 8'h00; 15'h4D21: d <= 8'h00; 15'h4D22: d <= 8'h00; 15'h4D23: d <= 8'h00;
                15'h4D24: d <= 8'h00; 15'h4D25: d <= 8'h00; 15'h4D26: d <= 8'h00; 15'h4D27: d <= 8'h00;
                15'h4D28: d <= 8'h00; 15'h4D29: d <= 8'h00; 15'h4D2A: d <= 8'h00; 15'h4D2B: d <= 8'h00;
                15'h4D2C: d <= 8'h00; 15'h4D2D: d <= 8'h00; 15'h4D2E: d <= 8'h00; 15'h4D2F: d <= 8'h7B;
                15'h4D30: d <= 8'h00; 15'h4D31: d <= 8'h00; 15'h4D32: d <= 8'h00; 15'h4D33: d <= 8'h00;
                15'h4D34: d <= 8'h00; 15'h4D35: d <= 8'h00; 15'h4D36: d <= 8'h00; 15'h4D37: d <= 8'h00;
                15'h4D38: d <= 8'h00; 15'h4D39: d <= 8'h00; 15'h4D3A: d <= 8'h00; 15'h4D3B: d <= 8'h00;
                15'h4D3C: d <= 8'h00; 15'h4D3D: d <= 8'h00; 15'h4D3E: d <= 8'h00; 15'h4D3F: d <= 8'h00;
                15'h4D40: d <= 8'h00; 15'h4D41: d <= 8'h00; 15'h4D42: d <= 8'h00; 15'h4D43: d <= 8'h00;
                15'h4D44: d <= 8'h00; 15'h4D45: d <= 8'h00; 15'h4D46: d <= 8'h00; 15'h4D47: d <= 8'h00;
                15'h4D48: d <= 8'h00; 15'h4D49: d <= 8'h00; 15'h4D4A: d <= 8'h00; 15'h4D4B: d <= 8'h00;
                15'h4D4C: d <= 8'h00; 15'h4D4D: d <= 8'h00; 15'h4D4E: d <= 8'h00; 15'h4D4F: d <= 8'h00;
                15'h4D50: d <= 8'h00; 15'h4D51: d <= 8'h00; 15'h4D52: d <= 8'h00; 15'h4D53: d <= 8'h00;
                15'h4D54: d <= 8'h00; 15'h4D55: d <= 8'h00; 15'h4D56: d <= 8'h00; 15'h4D57: d <= 8'h00;
                15'h4D58: d <= 8'h45; 15'h4D59: d <= 8'h35; 15'h4D5A: d <= 8'h32; 15'h4D5B: d <= 8'h00;
                15'h4D5C: d <= 8'h00; 15'h4D5D: d <= 8'h00; 15'h4D5E: d <= 8'h00; 15'h4D5F: d <= 8'h00;
                15'h4D60: d <= 8'h00; 15'h4D61: d <= 8'h00; 15'h4D62: d <= 8'h00; 15'h4D63: d <= 8'h00;
                15'h4D64: d <= 8'h00; 15'h4D65: d <= 8'h00; 15'h4D66: d <= 8'h00; 15'h4D67: d <= 8'h00;
                15'h4D68: d <= 8'h00; 15'h4D69: d <= 8'h00; 15'h4D6A: d <= 8'h00; 15'h4D6B: d <= 8'h00;
                15'h4D6C: d <= 8'h00; 15'h4D6D: d <= 8'h00; 15'h4D6E: d <= 8'h00; 15'h4D6F: d <= 8'h00;
                15'h4D70: d <= 8'h00; 15'h4D71: d <= 8'h00; 15'h4D72: d <= 8'h00; 15'h4D73: d <= 8'h00;
                15'h4D74: d <= 8'h00; 15'h4D75: d <= 8'h00; 15'h4D76: d <= 8'h00; 15'h4D77: d <= 8'h00;
                15'h4D78: d <= 8'h00; 15'h4D79: d <= 8'h00; 15'h4D7A: d <= 8'h00; 15'h4D7B: d <= 8'h00;
                15'h4D7C: d <= 8'h00; 15'h4D7D: d <= 8'h00; 15'h4D7E: d <= 8'h00; 15'h4D7F: d <= 8'hE0;
                15'h4D80: d <= 8'h10; 15'h4D81: d <= 8'h15; 15'h4D82: d <= 8'h1A; 15'h4D83: d <= 8'h1F;
                15'h4D84: d <= 8'h20; 15'h4D85: d <= 8'h25; 15'h4D86: d <= 8'h2A; 15'h4D87: d <= 8'h2F;
                15'h4D88: d <= 8'h34; 15'h4D89: d <= 8'h38; 15'h4D8A: d <= 8'h3C; 15'h4D8B: d <= 8'h31;
                15'h4D8C: d <= 8'h39; 15'h4D8D: d <= 8'h3D; 15'h4D8E: d <= 8'h32; 15'h4D8F: d <= 8'h36;
                15'h4D90: d <= 8'h3E; 15'h4D91: d <= 8'h33; 15'h4D92: d <= 8'h37; 15'h4D93: d <= 8'h3B;
                15'h4D94: d <= 8'h44; 15'h4D95: d <= 8'h48; 15'h4D96: d <= 8'h4C; 15'h4D97: d <= 8'h41;
                15'h4D98: d <= 8'h49; 15'h4D99: d <= 8'h4D; 15'h4D9A: d <= 8'h42; 15'h4D9B: d <= 8'h46;
                15'h4D9C: d <= 8'h4E; 15'h4D9D: d <= 8'h43; 15'h4D9E: d <= 8'h47; 15'h4D9F: d <= 8'h4B;
                15'h4DA0: d <= 8'h50; 15'h4DA1: d <= 8'h55; 15'h4DA2: d <= 8'h5A; 15'h4DA3: d <= 8'h5F;
                15'h4DA4: d <= 8'h60; 15'h4DA5: d <= 8'h65; 15'h4DA6: d <= 8'h6A; 15'h4DA7: d <= 8'h6F;
                15'h4DA8: d <= 8'h74; 15'h4DA9: d <= 8'h78; 15'h4DAA: d <= 8'h7C; 15'h4DAB: d <= 8'h71;
                15'h4DAC: d <= 8'h79; 15'h4DAD: d <= 8'h7D; 15'h4DAE: d <= 8'h72; 15'h4DAF: d <= 8'h76;
                15'h4DB0: d <= 8'h7E; 15'h4DB1: d <= 8'h73; 15'h4DB2: d <= 8'h77; 15'h4DB3: d <= 8'h7B;
                15'h4DB4: d <= 8'h84; 15'h4DB5: d <= 8'h88; 15'h4DB6: d <= 8'h8C; 15'h4DB7: d <= 8'h81;
                15'h4DB8: d <= 8'h89; 15'h4DB9: d <= 8'h8D; 15'h4DBA: d <= 8'h82; 15'h4DBB: d <= 8'h86;
                15'h4DBC: d <= 8'h8E; 15'h4DBD: d <= 8'h83; 15'h4DBE: d <= 8'h87; 15'h4DBF: d <= 8'h8B;
                15'h4DC0: d <= 8'h90; 15'h4DC1: d <= 8'h95; 15'h4DC2: d <= 8'h9A; 15'h4DC3: d <= 8'h9F;
                15'h4DC4: d <= 8'hA4; 15'h4DC5: d <= 8'hA8; 15'h4DC6: d <= 8'hAC; 15'h4DC7: d <= 8'hA1;
                15'h4DC8: d <= 8'hA9; 15'h4DC9: d <= 8'hAD; 15'h4DCA: d <= 8'hA2; 15'h4DCB: d <= 8'hA6;
                15'h4DCC: d <= 8'hAE; 15'h4DCD: d <= 8'hA3; 15'h4DCE: d <= 8'hA7; 15'h4DCF: d <= 8'hAB;
                15'h4DD0: d <= 8'hB4; 15'h4DD1: d <= 8'hB8; 15'h4DD2: d <= 8'hBC; 15'h4DD3: d <= 8'hB1;
                15'h4DD4: d <= 8'hB9; 15'h4DD5: d <= 8'hBD; 15'h4DD6: d <= 8'hB2; 15'h4DD7: d <= 8'hB6;
                15'h4DD8: d <= 8'hBE; 15'h4DD9: d <= 8'hB3; 15'h4DDA: d <= 8'hB7; 15'h4DDB: d <= 8'hBB;
                15'h4DDC: d <= 8'hC4; 15'h4DDD: d <= 8'hC8; 15'h4DDE: d <= 8'hCC; 15'h4DDF: d <= 8'hC1;
                15'h4DE0: d <= 8'hC9; 15'h4DE1: d <= 8'hCD; 15'h4DE2: d <= 8'hC2; 15'h4DE3: d <= 8'hC6;
                15'h4DE4: d <= 8'hCE; 15'h4DE5: d <= 8'hC3; 15'h4DE6: d <= 8'hC7; 15'h4DE7: d <= 8'hCB;
                15'h4DE8: d <= 8'hC0; 15'h4DE9: d <= 8'hC5; 15'h4DEA: d <= 8'hCA; 15'h4DEB: d <= 8'hCF;
                15'h4DEC: d <= 8'hD0; 15'h4DED: d <= 8'hD5; 15'h4DEE: d <= 8'hDA; 15'h4DEF: d <= 8'hDF;
                15'h4DF0: d <= 8'h74; 15'h4DF1: d <= 8'h78; 15'h4DF2: d <= 8'h7C; 15'h4DF3: d <= 8'h71;
                15'h4DF4: d <= 8'h79; 15'h4DF5: d <= 8'h7D; 15'h4DF6: d <= 8'h72; 15'h4DF7: d <= 8'h76;
                15'h4DF8: d <= 8'h7E; 15'h4DF9: d <= 8'h73; 15'h4DFA: d <= 8'h77; 15'h4DFB: d <= 8'h7B;
                15'h4DFC: d <= 8'hA0; 15'h4DFD: d <= 8'hA5; 15'h4DFE: d <= 8'hAA; 15'h4DFF: d <= 8'hAF;
                15'h4E00: d <= 8'h00; 15'h4E01: d <= 8'h00; 15'h4E02: d <= 8'h00; 15'h4E03: d <= 8'h00;
                15'h4E04: d <= 8'h00; 15'h4E05: d <= 8'h00; 15'h4E06: d <= 8'h00; 15'h4E07: d <= 8'h00;
                15'h4E08: d <= 8'h00; 15'h4E09: d <= 8'h00; 15'h4E0A: d <= 8'h00; 15'h4E0B: d <= 8'h00;
                15'h4E0C: d <= 8'h00; 15'h4E0D: d <= 8'h00; 15'h4E0E: d <= 8'h00; 15'h4E0F: d <= 8'h00;
                15'h4E10: d <= 8'h00; 15'h4E11: d <= 8'h00; 15'h4E12: d <= 8'h00; 15'h4E13: d <= 8'h00;
                15'h4E14: d <= 8'h00; 15'h4E15: d <= 8'h00; 15'h4E16: d <= 8'h00; 15'h4E17: d <= 8'h00;
                15'h4E18: d <= 8'h00; 15'h4E19: d <= 8'h00; 15'h4E1A: d <= 8'h00; 15'h4E1B: d <= 8'h00;
                15'h4E1C: d <= 8'h00; 15'h4E1D: d <= 8'h00; 15'h4E1E: d <= 8'h00; 15'h4E1F: d <= 8'h00;
                15'h4E20: d <= 8'h00; 15'h4E21: d <= 8'h00; 15'h4E22: d <= 8'h00; 15'h4E23: d <= 8'h00;
                15'h4E24: d <= 8'h00; 15'h4E25: d <= 8'h00; 15'h4E26: d <= 8'h00; 15'h4E27: d <= 8'h00;
                15'h4E28: d <= 8'h00; 15'h4E29: d <= 8'h00; 15'h4E2A: d <= 8'h00; 15'h4E2B: d <= 8'h00;
                15'h4E2C: d <= 8'h00; 15'h4E2D: d <= 8'h00; 15'h4E2E: d <= 8'h00; 15'h4E2F: d <= 8'h7B;
                15'h4E30: d <= 8'h00; 15'h4E31: d <= 8'h00; 15'h4E32: d <= 8'h00; 15'h4E33: d <= 8'h00;
                15'h4E34: d <= 8'h00; 15'h4E35: d <= 8'h00; 15'h4E36: d <= 8'h00; 15'h4E37: d <= 8'h00;
                15'h4E38: d <= 8'h00; 15'h4E39: d <= 8'h00; 15'h4E3A: d <= 8'h00; 15'h4E3B: d <= 8'h00;
                15'h4E3C: d <= 8'h00; 15'h4E3D: d <= 8'h00; 15'h4E3E: d <= 8'h00; 15'h4E3F: d <= 8'h00;
                15'h4E40: d <= 8'h00; 15'h4E41: d <= 8'h00; 15'h4E42: d <= 8'h00; 15'h4E43: d <= 8'h00;
                15'h4E44: d <= 8'h00; 15'h4E45: d <= 8'h00; 15'h4E46: d <= 8'h00; 15'h4E47: d <= 8'h00;
                15'h4E48: d <= 8'h00; 15'h4E49: d <= 8'h00; 15'h4E4A: d <= 8'h00; 15'h4E4B: d <= 8'h00;
                15'h4E4C: d <= 8'h00; 15'h4E4D: d <= 8'h00; 15'h4E4E: d <= 8'h00; 15'h4E4F: d <= 8'h00;
                15'h4E50: d <= 8'h00; 15'h4E51: d <= 8'h00; 15'h4E52: d <= 8'h00; 15'h4E53: d <= 8'h00;
                15'h4E54: d <= 8'h00; 15'h4E55: d <= 8'h00; 15'h4E56: d <= 8'h00; 15'h4E57: d <= 8'h00;
                15'h4E58: d <= 8'h45; 15'h4E59: d <= 8'h35; 15'h4E5A: d <= 8'h32; 15'h4E5B: d <= 8'h00;
                15'h4E5C: d <= 8'h00; 15'h4E5D: d <= 8'h00; 15'h4E5E: d <= 8'h00; 15'h4E5F: d <= 8'h00;
                15'h4E60: d <= 8'h00; 15'h4E61: d <= 8'h00; 15'h4E62: d <= 8'h00; 15'h4E63: d <= 8'h00;
                15'h4E64: d <= 8'h00; 15'h4E65: d <= 8'h00; 15'h4E66: d <= 8'h00; 15'h4E67: d <= 8'h00;
                15'h4E68: d <= 8'h00; 15'h4E69: d <= 8'h00; 15'h4E6A: d <= 8'h00; 15'h4E6B: d <= 8'h00;
                15'h4E6C: d <= 8'h00; 15'h4E6D: d <= 8'h00; 15'h4E6E: d <= 8'h00; 15'h4E6F: d <= 8'h00;
                15'h4E70: d <= 8'h00; 15'h4E71: d <= 8'h00; 15'h4E72: d <= 8'h00; 15'h4E73: d <= 8'h00;
                15'h4E74: d <= 8'h00; 15'h4E75: d <= 8'h00; 15'h4E76: d <= 8'h00; 15'h4E77: d <= 8'h00;
                15'h4E78: d <= 8'h00; 15'h4E79: d <= 8'h00; 15'h4E7A: d <= 8'h00; 15'h4E7B: d <= 8'h00;
                15'h4E7C: d <= 8'h00; 15'h4E7D: d <= 8'h00; 15'h4E7E: d <= 8'h00; 15'h4E7F: d <= 8'hE0;
                15'h4E80: d <= 8'h10; 15'h4E81: d <= 8'h15; 15'h4E82: d <= 8'h1A; 15'h4E83: d <= 8'h1F;
                15'h4E84: d <= 8'h20; 15'h4E85: d <= 8'h25; 15'h4E86: d <= 8'h2A; 15'h4E87: d <= 8'h2F;
                15'h4E88: d <= 8'h34; 15'h4E89: d <= 8'h38; 15'h4E8A: d <= 8'h3C; 15'h4E8B: d <= 8'h31;
                15'h4E8C: d <= 8'h39; 15'h4E8D: d <= 8'h3D; 15'h4E8E: d <= 8'h32; 15'h4E8F: d <= 8'h36;
                15'h4E90: d <= 8'h3E; 15'h4E91: d <= 8'h33; 15'h4E92: d <= 8'h37; 15'h4E93: d <= 8'h3B;
                15'h4E94: d <= 8'h44; 15'h4E95: d <= 8'h48; 15'h4E96: d <= 8'h4C; 15'h4E97: d <= 8'h41;
                15'h4E98: d <= 8'h49; 15'h4E99: d <= 8'h4D; 15'h4E9A: d <= 8'h42; 15'h4E9B: d <= 8'h46;
                15'h4E9C: d <= 8'h4E; 15'h4E9D: d <= 8'h43; 15'h4E9E: d <= 8'h47; 15'h4E9F: d <= 8'h4B;
                15'h4EA0: d <= 8'h50; 15'h4EA1: d <= 8'h55; 15'h4EA2: d <= 8'h5A; 15'h4EA3: d <= 8'h5F;
                15'h4EA4: d <= 8'h60; 15'h4EA5: d <= 8'h65; 15'h4EA6: d <= 8'h6A; 15'h4EA7: d <= 8'h6F;
                15'h4EA8: d <= 8'h74; 15'h4EA9: d <= 8'h78; 15'h4EAA: d <= 8'h7C; 15'h4EAB: d <= 8'h71;
                15'h4EAC: d <= 8'h79; 15'h4EAD: d <= 8'h7D; 15'h4EAE: d <= 8'h72; 15'h4EAF: d <= 8'h76;
                15'h4EB0: d <= 8'h7E; 15'h4EB1: d <= 8'h73; 15'h4EB2: d <= 8'h77; 15'h4EB3: d <= 8'h7B;
                15'h4EB4: d <= 8'h84; 15'h4EB5: d <= 8'h88; 15'h4EB6: d <= 8'h8C; 15'h4EB7: d <= 8'h81;
                15'h4EB8: d <= 8'h89; 15'h4EB9: d <= 8'h8D; 15'h4EBA: d <= 8'h82; 15'h4EBB: d <= 8'h86;
                15'h4EBC: d <= 8'h8E; 15'h4EBD: d <= 8'h83; 15'h4EBE: d <= 8'h87; 15'h4EBF: d <= 8'h8B;
                15'h4EC0: d <= 8'h90; 15'h4EC1: d <= 8'h95; 15'h4EC2: d <= 8'h9A; 15'h4EC3: d <= 8'h9F;
                15'h4EC4: d <= 8'hA4; 15'h4EC5: d <= 8'hA8; 15'h4EC6: d <= 8'hAC; 15'h4EC7: d <= 8'hA1;
                15'h4EC8: d <= 8'hA9; 15'h4EC9: d <= 8'hAD; 15'h4ECA: d <= 8'hA2; 15'h4ECB: d <= 8'hA6;
                15'h4ECC: d <= 8'hAE; 15'h4ECD: d <= 8'hA3; 15'h4ECE: d <= 8'hA7; 15'h4ECF: d <= 8'hAB;
                15'h4ED0: d <= 8'hB4; 15'h4ED1: d <= 8'hB8; 15'h4ED2: d <= 8'hBC; 15'h4ED3: d <= 8'hB1;
                15'h4ED4: d <= 8'hB9; 15'h4ED5: d <= 8'hBD; 15'h4ED6: d <= 8'hB2; 15'h4ED7: d <= 8'hB6;
                15'h4ED8: d <= 8'hBE; 15'h4ED9: d <= 8'hB3; 15'h4EDA: d <= 8'hB7; 15'h4EDB: d <= 8'hBB;
                15'h4EDC: d <= 8'hC4; 15'h4EDD: d <= 8'hC8; 15'h4EDE: d <= 8'hCC; 15'h4EDF: d <= 8'hC1;
                15'h4EE0: d <= 8'hC9; 15'h4EE1: d <= 8'hCD; 15'h4EE2: d <= 8'hC2; 15'h4EE3: d <= 8'hC6;
                15'h4EE4: d <= 8'hCE; 15'h4EE5: d <= 8'hC3; 15'h4EE6: d <= 8'hC7; 15'h4EE7: d <= 8'hCB;
                15'h4EE8: d <= 8'hC0; 15'h4EE9: d <= 8'hC5; 15'h4EEA: d <= 8'hCA; 15'h4EEB: d <= 8'hCF;
                15'h4EEC: d <= 8'hD0; 15'h4EED: d <= 8'hD5; 15'h4EEE: d <= 8'hDA; 15'h4EEF: d <= 8'hDF;
                15'h4EF0: d <= 8'h74; 15'h4EF1: d <= 8'h78; 15'h4EF2: d <= 8'h7C; 15'h4EF3: d <= 8'h71;
                15'h4EF4: d <= 8'h79; 15'h4EF5: d <= 8'h7D; 15'h4EF6: d <= 8'h72; 15'h4EF7: d <= 8'h76;
                15'h4EF8: d <= 8'h7E; 15'h4EF9: d <= 8'h73; 15'h4EFA: d <= 8'h77; 15'h4EFB: d <= 8'h7B;
                15'h4EFC: d <= 8'hA0; 15'h4EFD: d <= 8'hA5; 15'h4EFE: d <= 8'hAA; 15'h4EFF: d <= 8'hAF;
                15'h4F00: d <= 8'h00; 15'h4F01: d <= 8'h00; 15'h4F02: d <= 8'h00; 15'h4F03: d <= 8'h00;
                15'h4F04: d <= 8'h00; 15'h4F05: d <= 8'h00; 15'h4F06: d <= 8'h00; 15'h4F07: d <= 8'h00;
                15'h4F08: d <= 8'h00; 15'h4F09: d <= 8'h00; 15'h4F0A: d <= 8'h00; 15'h4F0B: d <= 8'h00;
                15'h4F0C: d <= 8'h00; 15'h4F0D: d <= 8'h00; 15'h4F0E: d <= 8'h00; 15'h4F0F: d <= 8'h00;
                15'h4F10: d <= 8'h00; 15'h4F11: d <= 8'h00; 15'h4F12: d <= 8'h00; 15'h4F13: d <= 8'h00;
                15'h4F14: d <= 8'h00; 15'h4F15: d <= 8'h00; 15'h4F16: d <= 8'h00; 15'h4F17: d <= 8'h00;
                15'h4F18: d <= 8'h00; 15'h4F19: d <= 8'h00; 15'h4F1A: d <= 8'h00; 15'h4F1B: d <= 8'h00;
                15'h4F1C: d <= 8'h00; 15'h4F1D: d <= 8'h00; 15'h4F1E: d <= 8'h00; 15'h4F1F: d <= 8'h00;
                15'h4F20: d <= 8'h00; 15'h4F21: d <= 8'h00; 15'h4F22: d <= 8'h00; 15'h4F23: d <= 8'h00;
                15'h4F24: d <= 8'h00; 15'h4F25: d <= 8'h00; 15'h4F26: d <= 8'h00; 15'h4F27: d <= 8'h00;
                15'h4F28: d <= 8'h00; 15'h4F29: d <= 8'h00; 15'h4F2A: d <= 8'h00; 15'h4F2B: d <= 8'h00;
                15'h4F2C: d <= 8'h00; 15'h4F2D: d <= 8'h00; 15'h4F2E: d <= 8'h00; 15'h4F2F: d <= 8'h7B;
                15'h4F30: d <= 8'h00; 15'h4F31: d <= 8'h00; 15'h4F32: d <= 8'h00; 15'h4F33: d <= 8'h00;
                15'h4F34: d <= 8'h00; 15'h4F35: d <= 8'h00; 15'h4F36: d <= 8'h00; 15'h4F37: d <= 8'h00;
                15'h4F38: d <= 8'h00; 15'h4F39: d <= 8'h00; 15'h4F3A: d <= 8'h00; 15'h4F3B: d <= 8'h00;
                15'h4F3C: d <= 8'h00; 15'h4F3D: d <= 8'h00; 15'h4F3E: d <= 8'h00; 15'h4F3F: d <= 8'h00;
                15'h4F40: d <= 8'h00; 15'h4F41: d <= 8'h00; 15'h4F42: d <= 8'h00; 15'h4F43: d <= 8'h00;
                15'h4F44: d <= 8'h00; 15'h4F45: d <= 8'h00; 15'h4F46: d <= 8'h00; 15'h4F47: d <= 8'h00;
                15'h4F48: d <= 8'h00; 15'h4F49: d <= 8'h00; 15'h4F4A: d <= 8'h00; 15'h4F4B: d <= 8'h00;
                15'h4F4C: d <= 8'h00; 15'h4F4D: d <= 8'h00; 15'h4F4E: d <= 8'h00; 15'h4F4F: d <= 8'h00;
                15'h4F50: d <= 8'h00; 15'h4F51: d <= 8'h00; 15'h4F52: d <= 8'h00; 15'h4F53: d <= 8'h00;
                15'h4F54: d <= 8'h00; 15'h4F55: d <= 8'h00; 15'h4F56: d <= 8'h00; 15'h4F57: d <= 8'h00;
                15'h4F58: d <= 8'h45; 15'h4F59: d <= 8'h35; 15'h4F5A: d <= 8'h32; 15'h4F5B: d <= 8'h00;
                15'h4F5C: d <= 8'h00; 15'h4F5D: d <= 8'h00; 15'h4F5E: d <= 8'h00; 15'h4F5F: d <= 8'h00;
                15'h4F60: d <= 8'h00; 15'h4F61: d <= 8'h00; 15'h4F62: d <= 8'h00; 15'h4F63: d <= 8'h00;
                15'h4F64: d <= 8'h00; 15'h4F65: d <= 8'h00; 15'h4F66: d <= 8'h00; 15'h4F67: d <= 8'h00;
                15'h4F68: d <= 8'h00; 15'h4F69: d <= 8'h00; 15'h4F6A: d <= 8'h00; 15'h4F6B: d <= 8'h00;
                15'h4F6C: d <= 8'h00; 15'h4F6D: d <= 8'h00; 15'h4F6E: d <= 8'h00; 15'h4F6F: d <= 8'h00;
                15'h4F70: d <= 8'h00; 15'h4F71: d <= 8'h00; 15'h4F72: d <= 8'h00; 15'h4F73: d <= 8'h00;
                15'h4F74: d <= 8'h00; 15'h4F75: d <= 8'h00; 15'h4F76: d <= 8'h00; 15'h4F77: d <= 8'h00;
                15'h4F78: d <= 8'h00; 15'h4F79: d <= 8'h00; 15'h4F7A: d <= 8'h00; 15'h4F7B: d <= 8'h00;
                15'h4F7C: d <= 8'h00; 15'h4F7D: d <= 8'h00; 15'h4F7E: d <= 8'h00; 15'h4F7F: d <= 8'hE0;
                15'h4F80: d <= 8'h10; 15'h4F81: d <= 8'h15; 15'h4F82: d <= 8'h1A; 15'h4F83: d <= 8'h1F;
                15'h4F84: d <= 8'h20; 15'h4F85: d <= 8'h25; 15'h4F86: d <= 8'h2A; 15'h4F87: d <= 8'h2F;
                15'h4F88: d <= 8'h34; 15'h4F89: d <= 8'h38; 15'h4F8A: d <= 8'h3C; 15'h4F8B: d <= 8'h31;
                15'h4F8C: d <= 8'h39; 15'h4F8D: d <= 8'h3D; 15'h4F8E: d <= 8'h32; 15'h4F8F: d <= 8'h36;
                15'h4F90: d <= 8'h3E; 15'h4F91: d <= 8'h33; 15'h4F92: d <= 8'h37; 15'h4F93: d <= 8'h3B;
                15'h4F94: d <= 8'h44; 15'h4F95: d <= 8'h48; 15'h4F96: d <= 8'h4C; 15'h4F97: d <= 8'h41;
                15'h4F98: d <= 8'h49; 15'h4F99: d <= 8'h4D; 15'h4F9A: d <= 8'h42; 15'h4F9B: d <= 8'h46;
                15'h4F9C: d <= 8'h4E; 15'h4F9D: d <= 8'h43; 15'h4F9E: d <= 8'h47; 15'h4F9F: d <= 8'h4B;
                15'h4FA0: d <= 8'h50; 15'h4FA1: d <= 8'h55; 15'h4FA2: d <= 8'h5A; 15'h4FA3: d <= 8'h5F;
                15'h4FA4: d <= 8'h60; 15'h4FA5: d <= 8'h65; 15'h4FA6: d <= 8'h6A; 15'h4FA7: d <= 8'h6F;
                15'h4FA8: d <= 8'h74; 15'h4FA9: d <= 8'h78; 15'h4FAA: d <= 8'h7C; 15'h4FAB: d <= 8'h71;
                15'h4FAC: d <= 8'h79; 15'h4FAD: d <= 8'h7D; 15'h4FAE: d <= 8'h72; 15'h4FAF: d <= 8'h76;
                15'h4FB0: d <= 8'h7E; 15'h4FB1: d <= 8'h73; 15'h4FB2: d <= 8'h77; 15'h4FB3: d <= 8'h7B;
                15'h4FB4: d <= 8'h84; 15'h4FB5: d <= 8'h88; 15'h4FB6: d <= 8'h8C; 15'h4FB7: d <= 8'h81;
                15'h4FB8: d <= 8'h89; 15'h4FB9: d <= 8'h8D; 15'h4FBA: d <= 8'h82; 15'h4FBB: d <= 8'h86;
                15'h4FBC: d <= 8'h8E; 15'h4FBD: d <= 8'h83; 15'h4FBE: d <= 8'h87; 15'h4FBF: d <= 8'h8B;
                15'h4FC0: d <= 8'h90; 15'h4FC1: d <= 8'h95; 15'h4FC2: d <= 8'h9A; 15'h4FC3: d <= 8'h9F;
                15'h4FC4: d <= 8'hA4; 15'h4FC5: d <= 8'hA8; 15'h4FC6: d <= 8'hAC; 15'h4FC7: d <= 8'hA1;
                15'h4FC8: d <= 8'hA9; 15'h4FC9: d <= 8'hAD; 15'h4FCA: d <= 8'hA2; 15'h4FCB: d <= 8'hA6;
                15'h4FCC: d <= 8'hAE; 15'h4FCD: d <= 8'hA3; 15'h4FCE: d <= 8'hA7; 15'h4FCF: d <= 8'hAB;
                15'h4FD0: d <= 8'hB4; 15'h4FD1: d <= 8'hB8; 15'h4FD2: d <= 8'hBC; 15'h4FD3: d <= 8'hB1;
                15'h4FD4: d <= 8'hB9; 15'h4FD5: d <= 8'hBD; 15'h4FD6: d <= 8'hB2; 15'h4FD7: d <= 8'hB6;
                15'h4FD8: d <= 8'hBE; 15'h4FD9: d <= 8'hB3; 15'h4FDA: d <= 8'hB7; 15'h4FDB: d <= 8'hBB;
                15'h4FDC: d <= 8'hC4; 15'h4FDD: d <= 8'hC8; 15'h4FDE: d <= 8'hCC; 15'h4FDF: d <= 8'hC1;
                15'h4FE0: d <= 8'hC9; 15'h4FE1: d <= 8'hCD; 15'h4FE2: d <= 8'hC2; 15'h4FE3: d <= 8'hC6;
                15'h4FE4: d <= 8'hCE; 15'h4FE5: d <= 8'hC3; 15'h4FE6: d <= 8'hC7; 15'h4FE7: d <= 8'hCB;
                15'h4FE8: d <= 8'hC0; 15'h4FE9: d <= 8'hC5; 15'h4FEA: d <= 8'hCA; 15'h4FEB: d <= 8'hCF;
                15'h4FEC: d <= 8'hD0; 15'h4FED: d <= 8'hD5; 15'h4FEE: d <= 8'hDA; 15'h4FEF: d <= 8'hDF;
                15'h4FF0: d <= 8'h74; 15'h4FF1: d <= 8'h78; 15'h4FF2: d <= 8'h7C; 15'h4FF3: d <= 8'h71;
                15'h4FF4: d <= 8'h79; 15'h4FF5: d <= 8'h7D; 15'h4FF6: d <= 8'h72; 15'h4FF7: d <= 8'h76;
                15'h4FF8: d <= 8'h7E; 15'h4FF9: d <= 8'h73; 15'h4FFA: d <= 8'h77; 15'h4FFB: d <= 8'h7B;
                15'h4FFC: d <= 8'hA0; 15'h4FFD: d <= 8'hA5; 15'h4FFE: d <= 8'hAA; 15'h4FFF: d <= 8'hAF;
                15'h5000: d <= 8'h00; 15'h5001: d <= 8'h00; 15'h5002: d <= 8'h00; 15'h5003: d <= 8'h00;
                15'h5004: d <= 8'h00; 15'h5005: d <= 8'h00; 15'h5006: d <= 8'h00; 15'h5007: d <= 8'h00;
                15'h5008: d <= 8'h00; 15'h5009: d <= 8'h00; 15'h500A: d <= 8'h00; 15'h500B: d <= 8'h00;
                15'h500C: d <= 8'h00; 15'h500D: d <= 8'h00; 15'h500E: d <= 8'h00; 15'h500F: d <= 8'h00;
                15'h5010: d <= 8'h00; 15'h5011: d <= 8'h00; 15'h5012: d <= 8'h00; 15'h5013: d <= 8'h00;
                15'h5014: d <= 8'h00; 15'h5015: d <= 8'h00; 15'h5016: d <= 8'h00; 15'h5017: d <= 8'h00;
                15'h5018: d <= 8'h00; 15'h5019: d <= 8'h00; 15'h501A: d <= 8'h00; 15'h501B: d <= 8'h00;
                15'h501C: d <= 8'h00; 15'h501D: d <= 8'h00; 15'h501E: d <= 8'h00; 15'h501F: d <= 8'h00;
                15'h5020: d <= 8'h00; 15'h5021: d <= 8'h00; 15'h5022: d <= 8'h00; 15'h5023: d <= 8'h00;
                15'h5024: d <= 8'h00; 15'h5025: d <= 8'h00; 15'h5026: d <= 8'h00; 15'h5027: d <= 8'h00;
                15'h5028: d <= 8'h00; 15'h5029: d <= 8'h00; 15'h502A: d <= 8'h00; 15'h502B: d <= 8'h00;
                15'h502C: d <= 8'h00; 15'h502D: d <= 8'h00; 15'h502E: d <= 8'h00; 15'h502F: d <= 8'hAF;
                15'h5030: d <= 8'h00; 15'h5031: d <= 8'h00; 15'h5032: d <= 8'h00; 15'h5033: d <= 8'h00;
                15'h5034: d <= 8'h00; 15'h5035: d <= 8'h00; 15'h5036: d <= 8'h00; 15'h5037: d <= 8'h00;
                15'h5038: d <= 8'h00; 15'h5039: d <= 8'h00; 15'h503A: d <= 8'h00; 15'h503B: d <= 8'h00;
                15'h503C: d <= 8'h00; 15'h503D: d <= 8'h00; 15'h503E: d <= 8'h00; 15'h503F: d <= 8'h00;
                15'h5040: d <= 8'h00; 15'h5041: d <= 8'h00; 15'h5042: d <= 8'h00; 15'h5043: d <= 8'h00;
                15'h5044: d <= 8'h00; 15'h5045: d <= 8'h00; 15'h5046: d <= 8'h00; 15'h5047: d <= 8'h00;
                15'h5048: d <= 8'h00; 15'h5049: d <= 8'h00; 15'h504A: d <= 8'h00; 15'h504B: d <= 8'h00;
                15'h504C: d <= 8'h00; 15'h504D: d <= 8'h00; 15'h504E: d <= 8'h00; 15'h504F: d <= 8'h00;
                15'h5050: d <= 8'h00; 15'h5051: d <= 8'h00; 15'h5052: d <= 8'h00; 15'h5053: d <= 8'h00;
                15'h5054: d <= 8'h00; 15'h5055: d <= 8'h00; 15'h5056: d <= 8'h00; 15'h5057: d <= 8'h00;
                15'h5058: d <= 8'h45; 15'h5059: d <= 8'h35; 15'h505A: d <= 8'hAA; 15'h505B: d <= 8'h00;
                15'h505C: d <= 8'h00; 15'h505D: d <= 8'h00; 15'h505E: d <= 8'h00; 15'h505F: d <= 8'h00;
                15'h5060: d <= 8'h00; 15'h5061: d <= 8'h00; 15'h5062: d <= 8'h00; 15'h5063: d <= 8'h00;
                15'h5064: d <= 8'h00; 15'h5065: d <= 8'h00; 15'h5066: d <= 8'h00; 15'h5067: d <= 8'h00;
                15'h5068: d <= 8'h00; 15'h5069: d <= 8'h00; 15'h506A: d <= 8'h00; 15'h506B: d <= 8'h00;
                15'h506C: d <= 8'h00; 15'h506D: d <= 8'h00; 15'h506E: d <= 8'h00; 15'h506F: d <= 8'h00;
                15'h5070: d <= 8'h00; 15'h5071: d <= 8'h00; 15'h5072: d <= 8'h00; 15'h5073: d <= 8'h00;
                15'h5074: d <= 8'h00; 15'h5075: d <= 8'h00; 15'h5076: d <= 8'h00; 15'h5077: d <= 8'h00;
                15'h5078: d <= 8'h00; 15'h5079: d <= 8'h00; 15'h507A: d <= 8'h00; 15'h507B: d <= 8'h00;
                15'h507C: d <= 8'h00; 15'h507D: d <= 8'h00; 15'h507E: d <= 8'h00; 15'h507F: d <= 8'hE0;
                15'h5080: d <= 8'h10; 15'h5081: d <= 8'h15; 15'h5082: d <= 8'h1A; 15'h5083: d <= 8'h1F;
                15'h5084: d <= 8'h20; 15'h5085: d <= 8'h25; 15'h5086: d <= 8'h2A; 15'h5087: d <= 8'h2F;
                15'h5088: d <= 8'h34; 15'h5089: d <= 8'h38; 15'h508A: d <= 8'h3C; 15'h508B: d <= 8'h31;
                15'h508C: d <= 8'h39; 15'h508D: d <= 8'h3D; 15'h508E: d <= 8'h32; 15'h508F: d <= 8'h36;
                15'h5090: d <= 8'h3E; 15'h5091: d <= 8'h33; 15'h5092: d <= 8'h37; 15'h5093: d <= 8'h3B;
                15'h5094: d <= 8'h44; 15'h5095: d <= 8'h48; 15'h5096: d <= 8'h4C; 15'h5097: d <= 8'h41;
                15'h5098: d <= 8'h49; 15'h5099: d <= 8'h4D; 15'h509A: d <= 8'h42; 15'h509B: d <= 8'h46;
                15'h509C: d <= 8'h4E; 15'h509D: d <= 8'h43; 15'h509E: d <= 8'h47; 15'h509F: d <= 8'h4B;
                15'h50A0: d <= 8'h50; 15'h50A1: d <= 8'h55; 15'h50A2: d <= 8'h5A; 15'h50A3: d <= 8'h5F;
                15'h50A4: d <= 8'h60; 15'h50A5: d <= 8'h65; 15'h50A6: d <= 8'h6A; 15'h50A7: d <= 8'h6F;
                15'h50A8: d <= 8'h74; 15'h50A9: d <= 8'h78; 15'h50AA: d <= 8'h7C; 15'h50AB: d <= 8'h71;
                15'h50AC: d <= 8'h79; 15'h50AD: d <= 8'h7D; 15'h50AE: d <= 8'h72; 15'h50AF: d <= 8'h76;
                15'h50B0: d <= 8'h7E; 15'h50B1: d <= 8'h73; 15'h50B2: d <= 8'h77; 15'h50B3: d <= 8'h7B;
                15'h50B4: d <= 8'h84; 15'h50B5: d <= 8'h88; 15'h50B6: d <= 8'h8C; 15'h50B7: d <= 8'h81;
                15'h50B8: d <= 8'h89; 15'h50B9: d <= 8'h8D; 15'h50BA: d <= 8'h82; 15'h50BB: d <= 8'h86;
                15'h50BC: d <= 8'h8E; 15'h50BD: d <= 8'h83; 15'h50BE: d <= 8'h87; 15'h50BF: d <= 8'h8B;
                15'h50C0: d <= 8'h90; 15'h50C1: d <= 8'h95; 15'h50C2: d <= 8'h9A; 15'h50C3: d <= 8'h9F;
                15'h50C4: d <= 8'hA4; 15'h50C5: d <= 8'hA8; 15'h50C6: d <= 8'hAC; 15'h50C7: d <= 8'hA1;
                15'h50C8: d <= 8'hA9; 15'h50C9: d <= 8'hAD; 15'h50CA: d <= 8'hA2; 15'h50CB: d <= 8'hA6;
                15'h50CC: d <= 8'hAE; 15'h50CD: d <= 8'hA3; 15'h50CE: d <= 8'hA7; 15'h50CF: d <= 8'hAB;
                15'h50D0: d <= 8'hB4; 15'h50D1: d <= 8'hB8; 15'h50D2: d <= 8'hBC; 15'h50D3: d <= 8'hB1;
                15'h50D4: d <= 8'hB9; 15'h50D5: d <= 8'hBD; 15'h50D6: d <= 8'hB2; 15'h50D7: d <= 8'hB6;
                15'h50D8: d <= 8'hBE; 15'h50D9: d <= 8'hB3; 15'h50DA: d <= 8'hB7; 15'h50DB: d <= 8'hBB;
                15'h50DC: d <= 8'hC4; 15'h50DD: d <= 8'hC8; 15'h50DE: d <= 8'hCC; 15'h50DF: d <= 8'hC1;
                15'h50E0: d <= 8'hC9; 15'h50E1: d <= 8'hCD; 15'h50E2: d <= 8'hC2; 15'h50E3: d <= 8'hC6;
                15'h50E4: d <= 8'hCE; 15'h50E5: d <= 8'hC3; 15'h50E6: d <= 8'hC7; 15'h50E7: d <= 8'hCB;
                15'h50E8: d <= 8'hC0; 15'h50E9: d <= 8'hC5; 15'h50EA: d <= 8'hCA; 15'h50EB: d <= 8'hCF;
                15'h50EC: d <= 8'hD0; 15'h50ED: d <= 8'hD5; 15'h50EE: d <= 8'hDA; 15'h50EF: d <= 8'hDF;
                15'h50F0: d <= 8'h74; 15'h50F1: d <= 8'h78; 15'h50F2: d <= 8'h7C; 15'h50F3: d <= 8'h71;
                15'h50F4: d <= 8'h79; 15'h50F5: d <= 8'h7D; 15'h50F6: d <= 8'h72; 15'h50F7: d <= 8'h76;
                15'h50F8: d <= 8'h7E; 15'h50F9: d <= 8'h73; 15'h50FA: d <= 8'h77; 15'h50FB: d <= 8'h7B;
                15'h50FC: d <= 8'hA0; 15'h50FD: d <= 8'hA5; 15'h50FE: d <= 8'hAA; 15'h50FF: d <= 8'hAF;
                15'h5100: d <= 8'h00; 15'h5101: d <= 8'h00; 15'h5102: d <= 8'h00; 15'h5103: d <= 8'h00;
                15'h5104: d <= 8'h00; 15'h5105: d <= 8'h00; 15'h5106: d <= 8'h00; 15'h5107: d <= 8'h00;
                15'h5108: d <= 8'h00; 15'h5109: d <= 8'h00; 15'h510A: d <= 8'h00; 15'h510B: d <= 8'h00;
                15'h510C: d <= 8'h00; 15'h510D: d <= 8'h00; 15'h510E: d <= 8'h00; 15'h510F: d <= 8'h00;
                15'h5110: d <= 8'h00; 15'h5111: d <= 8'h00; 15'h5112: d <= 8'h00; 15'h5113: d <= 8'h00;
                15'h5114: d <= 8'h00; 15'h5115: d <= 8'h00; 15'h5116: d <= 8'h00; 15'h5117: d <= 8'h00;
                15'h5118: d <= 8'h00; 15'h5119: d <= 8'h00; 15'h511A: d <= 8'h00; 15'h511B: d <= 8'h00;
                15'h511C: d <= 8'h00; 15'h511D: d <= 8'h00; 15'h511E: d <= 8'h00; 15'h511F: d <= 8'h00;
                15'h5120: d <= 8'h00; 15'h5121: d <= 8'h00; 15'h5122: d <= 8'h00; 15'h5123: d <= 8'h00;
                15'h5124: d <= 8'h00; 15'h5125: d <= 8'h00; 15'h5126: d <= 8'h00; 15'h5127: d <= 8'h00;
                15'h5128: d <= 8'h00; 15'h5129: d <= 8'h00; 15'h512A: d <= 8'h00; 15'h512B: d <= 8'h00;
                15'h512C: d <= 8'h00; 15'h512D: d <= 8'h00; 15'h512E: d <= 8'h00; 15'h512F: d <= 8'hAF;
                15'h5130: d <= 8'h00; 15'h5131: d <= 8'h00; 15'h5132: d <= 8'h00; 15'h5133: d <= 8'h00;
                15'h5134: d <= 8'h00; 15'h5135: d <= 8'h00; 15'h5136: d <= 8'h00; 15'h5137: d <= 8'h00;
                15'h5138: d <= 8'h00; 15'h5139: d <= 8'h00; 15'h513A: d <= 8'h00; 15'h513B: d <= 8'h00;
                15'h513C: d <= 8'h00; 15'h513D: d <= 8'h00; 15'h513E: d <= 8'h00; 15'h513F: d <= 8'h00;
                15'h5140: d <= 8'h00; 15'h5141: d <= 8'h00; 15'h5142: d <= 8'h00; 15'h5143: d <= 8'h00;
                15'h5144: d <= 8'h00; 15'h5145: d <= 8'h00; 15'h5146: d <= 8'h00; 15'h5147: d <= 8'h00;
                15'h5148: d <= 8'h00; 15'h5149: d <= 8'h00; 15'h514A: d <= 8'h00; 15'h514B: d <= 8'h00;
                15'h514C: d <= 8'h00; 15'h514D: d <= 8'h00; 15'h514E: d <= 8'h00; 15'h514F: d <= 8'h00;
                15'h5150: d <= 8'h00; 15'h5151: d <= 8'h00; 15'h5152: d <= 8'h00; 15'h5153: d <= 8'h00;
                15'h5154: d <= 8'h00; 15'h5155: d <= 8'h00; 15'h5156: d <= 8'h00; 15'h5157: d <= 8'h00;
                15'h5158: d <= 8'h45; 15'h5159: d <= 8'h35; 15'h515A: d <= 8'hAA; 15'h515B: d <= 8'h00;
                15'h515C: d <= 8'h00; 15'h515D: d <= 8'h00; 15'h515E: d <= 8'h00; 15'h515F: d <= 8'h00;
                15'h5160: d <= 8'h00; 15'h5161: d <= 8'h00; 15'h5162: d <= 8'h00; 15'h5163: d <= 8'h00;
                15'h5164: d <= 8'h00; 15'h5165: d <= 8'h00; 15'h5166: d <= 8'h00; 15'h5167: d <= 8'h00;
                15'h5168: d <= 8'h00; 15'h5169: d <= 8'h00; 15'h516A: d <= 8'h00; 15'h516B: d <= 8'h00;
                15'h516C: d <= 8'h00; 15'h516D: d <= 8'h00; 15'h516E: d <= 8'h00; 15'h516F: d <= 8'h00;
                15'h5170: d <= 8'h00; 15'h5171: d <= 8'h00; 15'h5172: d <= 8'h00; 15'h5173: d <= 8'h00;
                15'h5174: d <= 8'h00; 15'h5175: d <= 8'h00; 15'h5176: d <= 8'h00; 15'h5177: d <= 8'h00;
                15'h5178: d <= 8'h00; 15'h5179: d <= 8'h00; 15'h517A: d <= 8'h00; 15'h517B: d <= 8'h00;
                15'h517C: d <= 8'h00; 15'h517D: d <= 8'h00; 15'h517E: d <= 8'h00; 15'h517F: d <= 8'hE0;
                15'h5180: d <= 8'h10; 15'h5181: d <= 8'h15; 15'h5182: d <= 8'h1A; 15'h5183: d <= 8'h1F;
                15'h5184: d <= 8'h20; 15'h5185: d <= 8'h25; 15'h5186: d <= 8'h2A; 15'h5187: d <= 8'h2F;
                15'h5188: d <= 8'h34; 15'h5189: d <= 8'h38; 15'h518A: d <= 8'h3C; 15'h518B: d <= 8'h31;
                15'h518C: d <= 8'h39; 15'h518D: d <= 8'h3D; 15'h518E: d <= 8'h32; 15'h518F: d <= 8'h36;
                15'h5190: d <= 8'h3E; 15'h5191: d <= 8'h33; 15'h5192: d <= 8'h37; 15'h5193: d <= 8'h3B;
                15'h5194: d <= 8'h44; 15'h5195: d <= 8'h48; 15'h5196: d <= 8'h4C; 15'h5197: d <= 8'h41;
                15'h5198: d <= 8'h49; 15'h5199: d <= 8'h4D; 15'h519A: d <= 8'h42; 15'h519B: d <= 8'h46;
                15'h519C: d <= 8'h4E; 15'h519D: d <= 8'h43; 15'h519E: d <= 8'h47; 15'h519F: d <= 8'h4B;
                15'h51A0: d <= 8'h50; 15'h51A1: d <= 8'h55; 15'h51A2: d <= 8'h5A; 15'h51A3: d <= 8'h5F;
                15'h51A4: d <= 8'h60; 15'h51A5: d <= 8'h65; 15'h51A6: d <= 8'h6A; 15'h51A7: d <= 8'h6F;
                15'h51A8: d <= 8'h74; 15'h51A9: d <= 8'h78; 15'h51AA: d <= 8'h7C; 15'h51AB: d <= 8'h71;
                15'h51AC: d <= 8'h79; 15'h51AD: d <= 8'h7D; 15'h51AE: d <= 8'h72; 15'h51AF: d <= 8'h76;
                15'h51B0: d <= 8'h7E; 15'h51B1: d <= 8'h73; 15'h51B2: d <= 8'h77; 15'h51B3: d <= 8'h7B;
                15'h51B4: d <= 8'h84; 15'h51B5: d <= 8'h88; 15'h51B6: d <= 8'h8C; 15'h51B7: d <= 8'h81;
                15'h51B8: d <= 8'h89; 15'h51B9: d <= 8'h8D; 15'h51BA: d <= 8'h82; 15'h51BB: d <= 8'h86;
                15'h51BC: d <= 8'h8E; 15'h51BD: d <= 8'h83; 15'h51BE: d <= 8'h87; 15'h51BF: d <= 8'h8B;
                15'h51C0: d <= 8'h90; 15'h51C1: d <= 8'h95; 15'h51C2: d <= 8'h9A; 15'h51C3: d <= 8'h9F;
                15'h51C4: d <= 8'hA4; 15'h51C5: d <= 8'hA8; 15'h51C6: d <= 8'hAC; 15'h51C7: d <= 8'hA1;
                15'h51C8: d <= 8'hA9; 15'h51C9: d <= 8'hAD; 15'h51CA: d <= 8'hA2; 15'h51CB: d <= 8'hA6;
                15'h51CC: d <= 8'hAE; 15'h51CD: d <= 8'hA3; 15'h51CE: d <= 8'hA7; 15'h51CF: d <= 8'hAB;
                15'h51D0: d <= 8'hB4; 15'h51D1: d <= 8'hB8; 15'h51D2: d <= 8'hBC; 15'h51D3: d <= 8'hB1;
                15'h51D4: d <= 8'hB9; 15'h51D5: d <= 8'hBD; 15'h51D6: d <= 8'hB2; 15'h51D7: d <= 8'hB6;
                15'h51D8: d <= 8'hBE; 15'h51D9: d <= 8'hB3; 15'h51DA: d <= 8'hB7; 15'h51DB: d <= 8'hBB;
                15'h51DC: d <= 8'hC4; 15'h51DD: d <= 8'hC8; 15'h51DE: d <= 8'hCC; 15'h51DF: d <= 8'hC1;
                15'h51E0: d <= 8'hC9; 15'h51E1: d <= 8'hCD; 15'h51E2: d <= 8'hC2; 15'h51E3: d <= 8'hC6;
                15'h51E4: d <= 8'hCE; 15'h51E5: d <= 8'hC3; 15'h51E6: d <= 8'hC7; 15'h51E7: d <= 8'hCB;
                15'h51E8: d <= 8'hC0; 15'h51E9: d <= 8'hC5; 15'h51EA: d <= 8'hCA; 15'h51EB: d <= 8'hCF;
                15'h51EC: d <= 8'hD0; 15'h51ED: d <= 8'hD5; 15'h51EE: d <= 8'hDA; 15'h51EF: d <= 8'hDF;
                15'h51F0: d <= 8'h74; 15'h51F1: d <= 8'h78; 15'h51F2: d <= 8'h7C; 15'h51F3: d <= 8'h71;
                15'h51F4: d <= 8'h79; 15'h51F5: d <= 8'h7D; 15'h51F6: d <= 8'h72; 15'h51F7: d <= 8'h76;
                15'h51F8: d <= 8'h7E; 15'h51F9: d <= 8'h73; 15'h51FA: d <= 8'h77; 15'h51FB: d <= 8'h7B;
                15'h51FC: d <= 8'hA0; 15'h51FD: d <= 8'hA5; 15'h51FE: d <= 8'hAA; 15'h51FF: d <= 8'hAF;
                15'h5200: d <= 8'h00; 15'h5201: d <= 8'h00; 15'h5202: d <= 8'h00; 15'h5203: d <= 8'h00;
                15'h5204: d <= 8'h00; 15'h5205: d <= 8'h00; 15'h5206: d <= 8'h00; 15'h5207: d <= 8'h00;
                15'h5208: d <= 8'h00; 15'h5209: d <= 8'h00; 15'h520A: d <= 8'h00; 15'h520B: d <= 8'h00;
                15'h520C: d <= 8'h00; 15'h520D: d <= 8'h00; 15'h520E: d <= 8'h00; 15'h520F: d <= 8'h00;
                15'h5210: d <= 8'h00; 15'h5211: d <= 8'h00; 15'h5212: d <= 8'h00; 15'h5213: d <= 8'h00;
                15'h5214: d <= 8'h00; 15'h5215: d <= 8'h00; 15'h5216: d <= 8'h00; 15'h5217: d <= 8'h00;
                15'h5218: d <= 8'h00; 15'h5219: d <= 8'h00; 15'h521A: d <= 8'h00; 15'h521B: d <= 8'h00;
                15'h521C: d <= 8'h00; 15'h521D: d <= 8'h00; 15'h521E: d <= 8'h00; 15'h521F: d <= 8'h00;
                15'h5220: d <= 8'h00; 15'h5221: d <= 8'h00; 15'h5222: d <= 8'h00; 15'h5223: d <= 8'h00;
                15'h5224: d <= 8'h00; 15'h5225: d <= 8'h00; 15'h5226: d <= 8'h00; 15'h5227: d <= 8'h00;
                15'h5228: d <= 8'h00; 15'h5229: d <= 8'h00; 15'h522A: d <= 8'h00; 15'h522B: d <= 8'h00;
                15'h522C: d <= 8'h00; 15'h522D: d <= 8'h00; 15'h522E: d <= 8'h00; 15'h522F: d <= 8'hAF;
                15'h5230: d <= 8'h00; 15'h5231: d <= 8'h00; 15'h5232: d <= 8'h00; 15'h5233: d <= 8'h00;
                15'h5234: d <= 8'h00; 15'h5235: d <= 8'h00; 15'h5236: d <= 8'h00; 15'h5237: d <= 8'h00;
                15'h5238: d <= 8'h00; 15'h5239: d <= 8'h00; 15'h523A: d <= 8'h00; 15'h523B: d <= 8'h00;
                15'h523C: d <= 8'h00; 15'h523D: d <= 8'h00; 15'h523E: d <= 8'h00; 15'h523F: d <= 8'h00;
                15'h5240: d <= 8'h00; 15'h5241: d <= 8'h00; 15'h5242: d <= 8'h00; 15'h5243: d <= 8'h00;
                15'h5244: d <= 8'h00; 15'h5245: d <= 8'h00; 15'h5246: d <= 8'h00; 15'h5247: d <= 8'h00;
                15'h5248: d <= 8'h00; 15'h5249: d <= 8'h00; 15'h524A: d <= 8'h00; 15'h524B: d <= 8'h00;
                15'h524C: d <= 8'h00; 15'h524D: d <= 8'h00; 15'h524E: d <= 8'h00; 15'h524F: d <= 8'h00;
                15'h5250: d <= 8'h00; 15'h5251: d <= 8'h00; 15'h5252: d <= 8'h00; 15'h5253: d <= 8'h00;
                15'h5254: d <= 8'h00; 15'h5255: d <= 8'h00; 15'h5256: d <= 8'h00; 15'h5257: d <= 8'h00;
                15'h5258: d <= 8'h45; 15'h5259: d <= 8'h35; 15'h525A: d <= 8'hAA; 15'h525B: d <= 8'h00;
                15'h525C: d <= 8'h00; 15'h525D: d <= 8'h00; 15'h525E: d <= 8'h00; 15'h525F: d <= 8'h00;
                15'h5260: d <= 8'h00; 15'h5261: d <= 8'h00; 15'h5262: d <= 8'h00; 15'h5263: d <= 8'h00;
                15'h5264: d <= 8'h00; 15'h5265: d <= 8'h00; 15'h5266: d <= 8'h00; 15'h5267: d <= 8'h00;
                15'h5268: d <= 8'h00; 15'h5269: d <= 8'h00; 15'h526A: d <= 8'h00; 15'h526B: d <= 8'h00;
                15'h526C: d <= 8'h00; 15'h526D: d <= 8'h00; 15'h526E: d <= 8'h00; 15'h526F: d <= 8'h00;
                15'h5270: d <= 8'h00; 15'h5271: d <= 8'h00; 15'h5272: d <= 8'h00; 15'h5273: d <= 8'h00;
                15'h5274: d <= 8'h00; 15'h5275: d <= 8'h00; 15'h5276: d <= 8'h00; 15'h5277: d <= 8'h00;
                15'h5278: d <= 8'h00; 15'h5279: d <= 8'h00; 15'h527A: d <= 8'h00; 15'h527B: d <= 8'h00;
                15'h527C: d <= 8'h00; 15'h527D: d <= 8'h00; 15'h527E: d <= 8'h00; 15'h527F: d <= 8'hE0;
                15'h5280: d <= 8'h10; 15'h5281: d <= 8'h15; 15'h5282: d <= 8'h1A; 15'h5283: d <= 8'h1F;
                15'h5284: d <= 8'h20; 15'h5285: d <= 8'h25; 15'h5286: d <= 8'h2A; 15'h5287: d <= 8'h2F;
                15'h5288: d <= 8'h34; 15'h5289: d <= 8'h38; 15'h528A: d <= 8'h3C; 15'h528B: d <= 8'h31;
                15'h528C: d <= 8'h39; 15'h528D: d <= 8'h3D; 15'h528E: d <= 8'h32; 15'h528F: d <= 8'h36;
                15'h5290: d <= 8'h3E; 15'h5291: d <= 8'h33; 15'h5292: d <= 8'h37; 15'h5293: d <= 8'h3B;
                15'h5294: d <= 8'h44; 15'h5295: d <= 8'h48; 15'h5296: d <= 8'h4C; 15'h5297: d <= 8'h41;
                15'h5298: d <= 8'h49; 15'h5299: d <= 8'h4D; 15'h529A: d <= 8'h42; 15'h529B: d <= 8'h46;
                15'h529C: d <= 8'h4E; 15'h529D: d <= 8'h43; 15'h529E: d <= 8'h47; 15'h529F: d <= 8'h4B;
                15'h52A0: d <= 8'h50; 15'h52A1: d <= 8'h55; 15'h52A2: d <= 8'h5A; 15'h52A3: d <= 8'h5F;
                15'h52A4: d <= 8'h60; 15'h52A5: d <= 8'h65; 15'h52A6: d <= 8'h6A; 15'h52A7: d <= 8'h6F;
                15'h52A8: d <= 8'h74; 15'h52A9: d <= 8'h78; 15'h52AA: d <= 8'h7C; 15'h52AB: d <= 8'h71;
                15'h52AC: d <= 8'h79; 15'h52AD: d <= 8'h7D; 15'h52AE: d <= 8'h72; 15'h52AF: d <= 8'h76;
                15'h52B0: d <= 8'h7E; 15'h52B1: d <= 8'h73; 15'h52B2: d <= 8'h77; 15'h52B3: d <= 8'h7B;
                15'h52B4: d <= 8'h84; 15'h52B5: d <= 8'h88; 15'h52B6: d <= 8'h8C; 15'h52B7: d <= 8'h81;
                15'h52B8: d <= 8'h89; 15'h52B9: d <= 8'h8D; 15'h52BA: d <= 8'h82; 15'h52BB: d <= 8'h86;
                15'h52BC: d <= 8'h8E; 15'h52BD: d <= 8'h83; 15'h52BE: d <= 8'h87; 15'h52BF: d <= 8'h8B;
                15'h52C0: d <= 8'h90; 15'h52C1: d <= 8'h95; 15'h52C2: d <= 8'h9A; 15'h52C3: d <= 8'h9F;
                15'h52C4: d <= 8'hA4; 15'h52C5: d <= 8'hA8; 15'h52C6: d <= 8'hAC; 15'h52C7: d <= 8'hA1;
                15'h52C8: d <= 8'hA9; 15'h52C9: d <= 8'hAD; 15'h52CA: d <= 8'hA2; 15'h52CB: d <= 8'hA6;
                15'h52CC: d <= 8'hAE; 15'h52CD: d <= 8'hA3; 15'h52CE: d <= 8'hA7; 15'h52CF: d <= 8'hAB;
                15'h52D0: d <= 8'hB4; 15'h52D1: d <= 8'hB8; 15'h52D2: d <= 8'hBC; 15'h52D3: d <= 8'hB1;
                15'h52D4: d <= 8'hB9; 15'h52D5: d <= 8'hBD; 15'h52D6: d <= 8'hB2; 15'h52D7: d <= 8'hB6;
                15'h52D8: d <= 8'hBE; 15'h52D9: d <= 8'hB3; 15'h52DA: d <= 8'hB7; 15'h52DB: d <= 8'hBB;
                15'h52DC: d <= 8'hC4; 15'h52DD: d <= 8'hC8; 15'h52DE: d <= 8'hCC; 15'h52DF: d <= 8'hC1;
                15'h52E0: d <= 8'hC9; 15'h52E1: d <= 8'hCD; 15'h52E2: d <= 8'hC2; 15'h52E3: d <= 8'hC6;
                15'h52E4: d <= 8'hCE; 15'h52E5: d <= 8'hC3; 15'h52E6: d <= 8'hC7; 15'h52E7: d <= 8'hCB;
                15'h52E8: d <= 8'hC0; 15'h52E9: d <= 8'hC5; 15'h52EA: d <= 8'hCA; 15'h52EB: d <= 8'hCF;
                15'h52EC: d <= 8'hD0; 15'h52ED: d <= 8'hD5; 15'h52EE: d <= 8'hDA; 15'h52EF: d <= 8'hDF;
                15'h52F0: d <= 8'h74; 15'h52F1: d <= 8'h78; 15'h52F2: d <= 8'h7C; 15'h52F3: d <= 8'h71;
                15'h52F4: d <= 8'h79; 15'h52F5: d <= 8'h7D; 15'h52F6: d <= 8'h72; 15'h52F7: d <= 8'h76;
                15'h52F8: d <= 8'h7E; 15'h52F9: d <= 8'h73; 15'h52FA: d <= 8'h77; 15'h52FB: d <= 8'h7B;
                15'h52FC: d <= 8'hA0; 15'h52FD: d <= 8'hA5; 15'h52FE: d <= 8'hAA; 15'h52FF: d <= 8'hAF;
                15'h5300: d <= 8'h00; 15'h5301: d <= 8'h00; 15'h5302: d <= 8'h00; 15'h5303: d <= 8'h00;
                15'h5304: d <= 8'h00; 15'h5305: d <= 8'h00; 15'h5306: d <= 8'h00; 15'h5307: d <= 8'h00;
                15'h5308: d <= 8'h00; 15'h5309: d <= 8'h00; 15'h530A: d <= 8'h00; 15'h530B: d <= 8'h00;
                15'h530C: d <= 8'h00; 15'h530D: d <= 8'h00; 15'h530E: d <= 8'h00; 15'h530F: d <= 8'h00;
                15'h5310: d <= 8'h00; 15'h5311: d <= 8'h00; 15'h5312: d <= 8'h00; 15'h5313: d <= 8'h00;
                15'h5314: d <= 8'h00; 15'h5315: d <= 8'h00; 15'h5316: d <= 8'h00; 15'h5317: d <= 8'h00;
                15'h5318: d <= 8'h00; 15'h5319: d <= 8'h00; 15'h531A: d <= 8'h00; 15'h531B: d <= 8'h00;
                15'h531C: d <= 8'h00; 15'h531D: d <= 8'h00; 15'h531E: d <= 8'h00; 15'h531F: d <= 8'h00;
                15'h5320: d <= 8'h00; 15'h5321: d <= 8'h00; 15'h5322: d <= 8'h00; 15'h5323: d <= 8'h00;
                15'h5324: d <= 8'h00; 15'h5325: d <= 8'h00; 15'h5326: d <= 8'h00; 15'h5327: d <= 8'h00;
                15'h5328: d <= 8'h00; 15'h5329: d <= 8'h00; 15'h532A: d <= 8'h00; 15'h532B: d <= 8'h00;
                15'h532C: d <= 8'h00; 15'h532D: d <= 8'h00; 15'h532E: d <= 8'h00; 15'h532F: d <= 8'hAF;
                15'h5330: d <= 8'h00; 15'h5331: d <= 8'h00; 15'h5332: d <= 8'h00; 15'h5333: d <= 8'h00;
                15'h5334: d <= 8'h00; 15'h5335: d <= 8'h00; 15'h5336: d <= 8'h00; 15'h5337: d <= 8'h00;
                15'h5338: d <= 8'h00; 15'h5339: d <= 8'h00; 15'h533A: d <= 8'h00; 15'h533B: d <= 8'h00;
                15'h533C: d <= 8'h00; 15'h533D: d <= 8'h00; 15'h533E: d <= 8'h00; 15'h533F: d <= 8'h00;
                15'h5340: d <= 8'h00; 15'h5341: d <= 8'h00; 15'h5342: d <= 8'h00; 15'h5343: d <= 8'h00;
                15'h5344: d <= 8'h00; 15'h5345: d <= 8'h00; 15'h5346: d <= 8'h00; 15'h5347: d <= 8'h00;
                15'h5348: d <= 8'h00; 15'h5349: d <= 8'h00; 15'h534A: d <= 8'h00; 15'h534B: d <= 8'h00;
                15'h534C: d <= 8'h00; 15'h534D: d <= 8'h00; 15'h534E: d <= 8'h00; 15'h534F: d <= 8'h00;
                15'h5350: d <= 8'h00; 15'h5351: d <= 8'h00; 15'h5352: d <= 8'h00; 15'h5353: d <= 8'h00;
                15'h5354: d <= 8'h00; 15'h5355: d <= 8'h00; 15'h5356: d <= 8'h00; 15'h5357: d <= 8'h00;
                15'h5358: d <= 8'h45; 15'h5359: d <= 8'h35; 15'h535A: d <= 8'hAA; 15'h535B: d <= 8'h00;
                15'h535C: d <= 8'h00; 15'h535D: d <= 8'h00; 15'h535E: d <= 8'h00; 15'h535F: d <= 8'h00;
                15'h5360: d <= 8'h00; 15'h5361: d <= 8'h00; 15'h5362: d <= 8'h00; 15'h5363: d <= 8'h00;
                15'h5364: d <= 8'h00; 15'h5365: d <= 8'h00; 15'h5366: d <= 8'h00; 15'h5367: d <= 8'h00;
                15'h5368: d <= 8'h00; 15'h5369: d <= 8'h00; 15'h536A: d <= 8'h00; 15'h536B: d <= 8'h00;
                15'h536C: d <= 8'h00; 15'h536D: d <= 8'h00; 15'h536E: d <= 8'h00; 15'h536F: d <= 8'h00;
                15'h5370: d <= 8'h00; 15'h5371: d <= 8'h00; 15'h5372: d <= 8'h00; 15'h5373: d <= 8'h00;
                15'h5374: d <= 8'h00; 15'h5375: d <= 8'h00; 15'h5376: d <= 8'h00; 15'h5377: d <= 8'h00;
                15'h5378: d <= 8'h00; 15'h5379: d <= 8'h00; 15'h537A: d <= 8'h00; 15'h537B: d <= 8'h00;
                15'h537C: d <= 8'h00; 15'h537D: d <= 8'h00; 15'h537E: d <= 8'h00; 15'h537F: d <= 8'hE0;
                15'h5380: d <= 8'h10; 15'h5381: d <= 8'h15; 15'h5382: d <= 8'h1A; 15'h5383: d <= 8'h1F;
                15'h5384: d <= 8'h20; 15'h5385: d <= 8'h25; 15'h5386: d <= 8'h2A; 15'h5387: d <= 8'h2F;
                15'h5388: d <= 8'h34; 15'h5389: d <= 8'h38; 15'h538A: d <= 8'h3C; 15'h538B: d <= 8'h31;
                15'h538C: d <= 8'h39; 15'h538D: d <= 8'h3D; 15'h538E: d <= 8'h32; 15'h538F: d <= 8'h36;
                15'h5390: d <= 8'h3E; 15'h5391: d <= 8'h33; 15'h5392: d <= 8'h37; 15'h5393: d <= 8'h3B;
                15'h5394: d <= 8'h44; 15'h5395: d <= 8'h48; 15'h5396: d <= 8'h4C; 15'h5397: d <= 8'h41;
                15'h5398: d <= 8'h49; 15'h5399: d <= 8'h4D; 15'h539A: d <= 8'h42; 15'h539B: d <= 8'h46;
                15'h539C: d <= 8'h4E; 15'h539D: d <= 8'h43; 15'h539E: d <= 8'h47; 15'h539F: d <= 8'h4B;
                15'h53A0: d <= 8'h50; 15'h53A1: d <= 8'h55; 15'h53A2: d <= 8'h5A; 15'h53A3: d <= 8'h5F;
                15'h53A4: d <= 8'h60; 15'h53A5: d <= 8'h65; 15'h53A6: d <= 8'h6A; 15'h53A7: d <= 8'h6F;
                15'h53A8: d <= 8'h74; 15'h53A9: d <= 8'h78; 15'h53AA: d <= 8'h7C; 15'h53AB: d <= 8'h71;
                15'h53AC: d <= 8'h79; 15'h53AD: d <= 8'h7D; 15'h53AE: d <= 8'h72; 15'h53AF: d <= 8'h76;
                15'h53B0: d <= 8'h7E; 15'h53B1: d <= 8'h73; 15'h53B2: d <= 8'h77; 15'h53B3: d <= 8'h7B;
                15'h53B4: d <= 8'h84; 15'h53B5: d <= 8'h88; 15'h53B6: d <= 8'h8C; 15'h53B7: d <= 8'h81;
                15'h53B8: d <= 8'h89; 15'h53B9: d <= 8'h8D; 15'h53BA: d <= 8'h82; 15'h53BB: d <= 8'h86;
                15'h53BC: d <= 8'h8E; 15'h53BD: d <= 8'h83; 15'h53BE: d <= 8'h87; 15'h53BF: d <= 8'h8B;
                15'h53C0: d <= 8'h90; 15'h53C1: d <= 8'h95; 15'h53C2: d <= 8'h9A; 15'h53C3: d <= 8'h9F;
                15'h53C4: d <= 8'hA4; 15'h53C5: d <= 8'hA8; 15'h53C6: d <= 8'hAC; 15'h53C7: d <= 8'hA1;
                15'h53C8: d <= 8'hA9; 15'h53C9: d <= 8'hAD; 15'h53CA: d <= 8'hA2; 15'h53CB: d <= 8'hA6;
                15'h53CC: d <= 8'hAE; 15'h53CD: d <= 8'hA3; 15'h53CE: d <= 8'hA7; 15'h53CF: d <= 8'hAB;
                15'h53D0: d <= 8'hB4; 15'h53D1: d <= 8'hB8; 15'h53D2: d <= 8'hBC; 15'h53D3: d <= 8'hB1;
                15'h53D4: d <= 8'hB9; 15'h53D5: d <= 8'hBD; 15'h53D6: d <= 8'hB2; 15'h53D7: d <= 8'hB6;
                15'h53D8: d <= 8'hBE; 15'h53D9: d <= 8'hB3; 15'h53DA: d <= 8'hB7; 15'h53DB: d <= 8'hBB;
                15'h53DC: d <= 8'hC4; 15'h53DD: d <= 8'hC8; 15'h53DE: d <= 8'hCC; 15'h53DF: d <= 8'hC1;
                15'h53E0: d <= 8'hC9; 15'h53E1: d <= 8'hCD; 15'h53E2: d <= 8'hC2; 15'h53E3: d <= 8'hC6;
                15'h53E4: d <= 8'hCE; 15'h53E5: d <= 8'hC3; 15'h53E6: d <= 8'hC7; 15'h53E7: d <= 8'hCB;
                15'h53E8: d <= 8'hC0; 15'h53E9: d <= 8'hC5; 15'h53EA: d <= 8'hCA; 15'h53EB: d <= 8'hCF;
                15'h53EC: d <= 8'hD0; 15'h53ED: d <= 8'hD5; 15'h53EE: d <= 8'hDA; 15'h53EF: d <= 8'hDF;
                15'h53F0: d <= 8'h74; 15'h53F1: d <= 8'h78; 15'h53F2: d <= 8'h7C; 15'h53F3: d <= 8'h71;
                15'h53F4: d <= 8'h79; 15'h53F5: d <= 8'h7D; 15'h53F6: d <= 8'h72; 15'h53F7: d <= 8'h76;
                15'h53F8: d <= 8'h7E; 15'h53F9: d <= 8'h73; 15'h53FA: d <= 8'h77; 15'h53FB: d <= 8'h7B;
                15'h53FC: d <= 8'hA0; 15'h53FD: d <= 8'hA5; 15'h53FE: d <= 8'hAA; 15'h53FF: d <= 8'hAF;
                15'h5400: d <= 8'h00; 15'h5401: d <= 8'h00; 15'h5402: d <= 8'h00; 15'h5403: d <= 8'h00;
                15'h5404: d <= 8'h00; 15'h5405: d <= 8'h00; 15'h5406: d <= 8'h00; 15'h5407: d <= 8'h00;
                15'h5408: d <= 8'h00; 15'h5409: d <= 8'h00; 15'h540A: d <= 8'h00; 15'h540B: d <= 8'h00;
                15'h540C: d <= 8'h00; 15'h540D: d <= 8'h00; 15'h540E: d <= 8'h00; 15'h540F: d <= 8'h00;
                15'h5410: d <= 8'h00; 15'h5411: d <= 8'h00; 15'h5412: d <= 8'h00; 15'h5413: d <= 8'h00;
                15'h5414: d <= 8'h00; 15'h5415: d <= 8'h00; 15'h5416: d <= 8'h00; 15'h5417: d <= 8'h00;
                15'h5418: d <= 8'h00; 15'h5419: d <= 8'h00; 15'h541A: d <= 8'h00; 15'h541B: d <= 8'h00;
                15'h541C: d <= 8'h00; 15'h541D: d <= 8'h00; 15'h541E: d <= 8'h00; 15'h541F: d <= 8'h00;
                15'h5420: d <= 8'h00; 15'h5421: d <= 8'h00; 15'h5422: d <= 8'h00; 15'h5423: d <= 8'h00;
                15'h5424: d <= 8'h00; 15'h5425: d <= 8'h00; 15'h5426: d <= 8'h00; 15'h5427: d <= 8'h00;
                15'h5428: d <= 8'h00; 15'h5429: d <= 8'h00; 15'h542A: d <= 8'h00; 15'h542B: d <= 8'h00;
                15'h542C: d <= 8'h00; 15'h542D: d <= 8'h00; 15'h542E: d <= 8'h00; 15'h542F: d <= 8'hAF;
                15'h5430: d <= 8'h00; 15'h5431: d <= 8'h00; 15'h5432: d <= 8'h00; 15'h5433: d <= 8'h00;
                15'h5434: d <= 8'h00; 15'h5435: d <= 8'h00; 15'h5436: d <= 8'h00; 15'h5437: d <= 8'h00;
                15'h5438: d <= 8'h00; 15'h5439: d <= 8'h00; 15'h543A: d <= 8'h00; 15'h543B: d <= 8'h00;
                15'h543C: d <= 8'h00; 15'h543D: d <= 8'h00; 15'h543E: d <= 8'h00; 15'h543F: d <= 8'h00;
                15'h5440: d <= 8'h00; 15'h5441: d <= 8'h00; 15'h5442: d <= 8'h00; 15'h5443: d <= 8'h00;
                15'h5444: d <= 8'h00; 15'h5445: d <= 8'h00; 15'h5446: d <= 8'h00; 15'h5447: d <= 8'h00;
                15'h5448: d <= 8'h00; 15'h5449: d <= 8'h00; 15'h544A: d <= 8'h00; 15'h544B: d <= 8'h00;
                15'h544C: d <= 8'h00; 15'h544D: d <= 8'h00; 15'h544E: d <= 8'h00; 15'h544F: d <= 8'h00;
                15'h5450: d <= 8'h00; 15'h5451: d <= 8'h00; 15'h5452: d <= 8'h00; 15'h5453: d <= 8'h00;
                15'h5454: d <= 8'h00; 15'h5455: d <= 8'h00; 15'h5456: d <= 8'h00; 15'h5457: d <= 8'h00;
                15'h5458: d <= 8'h45; 15'h5459: d <= 8'h35; 15'h545A: d <= 8'hAA; 15'h545B: d <= 8'h00;
                15'h545C: d <= 8'h00; 15'h545D: d <= 8'h00; 15'h545E: d <= 8'h00; 15'h545F: d <= 8'h00;
                15'h5460: d <= 8'h00; 15'h5461: d <= 8'h00; 15'h5462: d <= 8'h00; 15'h5463: d <= 8'h00;
                15'h5464: d <= 8'h00; 15'h5465: d <= 8'h00; 15'h5466: d <= 8'h00; 15'h5467: d <= 8'h00;
                15'h5468: d <= 8'h00; 15'h5469: d <= 8'h00; 15'h546A: d <= 8'h00; 15'h546B: d <= 8'h00;
                15'h546C: d <= 8'h00; 15'h546D: d <= 8'h00; 15'h546E: d <= 8'h00; 15'h546F: d <= 8'h00;
                15'h5470: d <= 8'h00; 15'h5471: d <= 8'h00; 15'h5472: d <= 8'h00; 15'h5473: d <= 8'h00;
                15'h5474: d <= 8'h00; 15'h5475: d <= 8'h00; 15'h5476: d <= 8'h00; 15'h5477: d <= 8'h00;
                15'h5478: d <= 8'h00; 15'h5479: d <= 8'h00; 15'h547A: d <= 8'h00; 15'h547B: d <= 8'h00;
                15'h547C: d <= 8'h00; 15'h547D: d <= 8'h00; 15'h547E: d <= 8'h00; 15'h547F: d <= 8'hE0;
                15'h5480: d <= 8'h10; 15'h5481: d <= 8'h15; 15'h5482: d <= 8'h1A; 15'h5483: d <= 8'h1F;
                15'h5484: d <= 8'h20; 15'h5485: d <= 8'h25; 15'h5486: d <= 8'h2A; 15'h5487: d <= 8'h2F;
                15'h5488: d <= 8'h34; 15'h5489: d <= 8'h38; 15'h548A: d <= 8'h3C; 15'h548B: d <= 8'h31;
                15'h548C: d <= 8'h39; 15'h548D: d <= 8'h3D; 15'h548E: d <= 8'h32; 15'h548F: d <= 8'h36;
                15'h5490: d <= 8'h3E; 15'h5491: d <= 8'h33; 15'h5492: d <= 8'h37; 15'h5493: d <= 8'h3B;
                15'h5494: d <= 8'h44; 15'h5495: d <= 8'h48; 15'h5496: d <= 8'h4C; 15'h5497: d <= 8'h41;
                15'h5498: d <= 8'h49; 15'h5499: d <= 8'h4D; 15'h549A: d <= 8'h42; 15'h549B: d <= 8'h46;
                15'h549C: d <= 8'h4E; 15'h549D: d <= 8'h43; 15'h549E: d <= 8'h47; 15'h549F: d <= 8'h4B;
                15'h54A0: d <= 8'h50; 15'h54A1: d <= 8'h55; 15'h54A2: d <= 8'h5A; 15'h54A3: d <= 8'h5F;
                15'h54A4: d <= 8'h60; 15'h54A5: d <= 8'h65; 15'h54A6: d <= 8'h6A; 15'h54A7: d <= 8'h6F;
                15'h54A8: d <= 8'h74; 15'h54A9: d <= 8'h78; 15'h54AA: d <= 8'h7C; 15'h54AB: d <= 8'h71;
                15'h54AC: d <= 8'h79; 15'h54AD: d <= 8'h7D; 15'h54AE: d <= 8'h72; 15'h54AF: d <= 8'h76;
                15'h54B0: d <= 8'h7E; 15'h54B1: d <= 8'h73; 15'h54B2: d <= 8'h77; 15'h54B3: d <= 8'h7B;
                15'h54B4: d <= 8'h84; 15'h54B5: d <= 8'h88; 15'h54B6: d <= 8'h8C; 15'h54B7: d <= 8'h81;
                15'h54B8: d <= 8'h89; 15'h54B9: d <= 8'h8D; 15'h54BA: d <= 8'h82; 15'h54BB: d <= 8'h86;
                15'h54BC: d <= 8'h8E; 15'h54BD: d <= 8'h83; 15'h54BE: d <= 8'h87; 15'h54BF: d <= 8'h8B;
                15'h54C0: d <= 8'h90; 15'h54C1: d <= 8'h95; 15'h54C2: d <= 8'h9A; 15'h54C3: d <= 8'h9F;
                15'h54C4: d <= 8'hA4; 15'h54C5: d <= 8'hA8; 15'h54C6: d <= 8'hAC; 15'h54C7: d <= 8'hA1;
                15'h54C8: d <= 8'hA9; 15'h54C9: d <= 8'hAD; 15'h54CA: d <= 8'hA2; 15'h54CB: d <= 8'hA6;
                15'h54CC: d <= 8'hAE; 15'h54CD: d <= 8'hA3; 15'h54CE: d <= 8'hA7; 15'h54CF: d <= 8'hAB;
                15'h54D0: d <= 8'hB4; 15'h54D1: d <= 8'hB8; 15'h54D2: d <= 8'hBC; 15'h54D3: d <= 8'hB1;
                15'h54D4: d <= 8'hB9; 15'h54D5: d <= 8'hBD; 15'h54D6: d <= 8'hB2; 15'h54D7: d <= 8'hB6;
                15'h54D8: d <= 8'hBE; 15'h54D9: d <= 8'hB3; 15'h54DA: d <= 8'hB7; 15'h54DB: d <= 8'hBB;
                15'h54DC: d <= 8'hC4; 15'h54DD: d <= 8'hC8; 15'h54DE: d <= 8'hCC; 15'h54DF: d <= 8'hC1;
                15'h54E0: d <= 8'hC9; 15'h54E1: d <= 8'hCD; 15'h54E2: d <= 8'hC2; 15'h54E3: d <= 8'hC6;
                15'h54E4: d <= 8'hCE; 15'h54E5: d <= 8'hC3; 15'h54E6: d <= 8'hC7; 15'h54E7: d <= 8'hCB;
                15'h54E8: d <= 8'hC0; 15'h54E9: d <= 8'hC5; 15'h54EA: d <= 8'hCA; 15'h54EB: d <= 8'hCF;
                15'h54EC: d <= 8'hD0; 15'h54ED: d <= 8'hD5; 15'h54EE: d <= 8'hDA; 15'h54EF: d <= 8'hDF;
                15'h54F0: d <= 8'h74; 15'h54F1: d <= 8'h78; 15'h54F2: d <= 8'h7C; 15'h54F3: d <= 8'h71;
                15'h54F4: d <= 8'h79; 15'h54F5: d <= 8'h7D; 15'h54F6: d <= 8'h72; 15'h54F7: d <= 8'h76;
                15'h54F8: d <= 8'h7E; 15'h54F9: d <= 8'h73; 15'h54FA: d <= 8'h77; 15'h54FB: d <= 8'h7B;
                15'h54FC: d <= 8'hA0; 15'h54FD: d <= 8'hA5; 15'h54FE: d <= 8'hAA; 15'h54FF: d <= 8'hAF;
                15'h5500: d <= 8'h00; 15'h5501: d <= 8'h00; 15'h5502: d <= 8'h00; 15'h5503: d <= 8'h00;
                15'h5504: d <= 8'h00; 15'h5505: d <= 8'h00; 15'h5506: d <= 8'h00; 15'h5507: d <= 8'h00;
                15'h5508: d <= 8'h00; 15'h5509: d <= 8'h00; 15'h550A: d <= 8'h00; 15'h550B: d <= 8'h00;
                15'h550C: d <= 8'h00; 15'h550D: d <= 8'h00; 15'h550E: d <= 8'h00; 15'h550F: d <= 8'h00;
                15'h5510: d <= 8'h00; 15'h5511: d <= 8'h00; 15'h5512: d <= 8'h00; 15'h5513: d <= 8'h00;
                15'h5514: d <= 8'h00; 15'h5515: d <= 8'h00; 15'h5516: d <= 8'h00; 15'h5517: d <= 8'h00;
                15'h5518: d <= 8'h00; 15'h5519: d <= 8'h00; 15'h551A: d <= 8'h00; 15'h551B: d <= 8'h00;
                15'h551C: d <= 8'h00; 15'h551D: d <= 8'h00; 15'h551E: d <= 8'h00; 15'h551F: d <= 8'h00;
                15'h5520: d <= 8'h00; 15'h5521: d <= 8'h00; 15'h5522: d <= 8'h00; 15'h5523: d <= 8'h00;
                15'h5524: d <= 8'h00; 15'h5525: d <= 8'h00; 15'h5526: d <= 8'h00; 15'h5527: d <= 8'h00;
                15'h5528: d <= 8'h00; 15'h5529: d <= 8'h00; 15'h552A: d <= 8'h00; 15'h552B: d <= 8'h00;
                15'h552C: d <= 8'h00; 15'h552D: d <= 8'h00; 15'h552E: d <= 8'h00; 15'h552F: d <= 8'hAF;
                15'h5530: d <= 8'h00; 15'h5531: d <= 8'h00; 15'h5532: d <= 8'h00; 15'h5533: d <= 8'h00;
                15'h5534: d <= 8'h00; 15'h5535: d <= 8'h00; 15'h5536: d <= 8'h00; 15'h5537: d <= 8'h00;
                15'h5538: d <= 8'h00; 15'h5539: d <= 8'h00; 15'h553A: d <= 8'h00; 15'h553B: d <= 8'h00;
                15'h553C: d <= 8'h00; 15'h553D: d <= 8'h00; 15'h553E: d <= 8'h00; 15'h553F: d <= 8'h00;
                15'h5540: d <= 8'h00; 15'h5541: d <= 8'h00; 15'h5542: d <= 8'h00; 15'h5543: d <= 8'h00;
                15'h5544: d <= 8'h00; 15'h5545: d <= 8'h00; 15'h5546: d <= 8'h00; 15'h5547: d <= 8'h00;
                15'h5548: d <= 8'h00; 15'h5549: d <= 8'h00; 15'h554A: d <= 8'h00; 15'h554B: d <= 8'h00;
                15'h554C: d <= 8'h00; 15'h554D: d <= 8'h00; 15'h554E: d <= 8'h00; 15'h554F: d <= 8'h00;
                15'h5550: d <= 8'h00; 15'h5551: d <= 8'h00; 15'h5552: d <= 8'h00; 15'h5553: d <= 8'h00;
                15'h5554: d <= 8'h00; 15'h5555: d <= 8'h00; 15'h5556: d <= 8'h00; 15'h5557: d <= 8'h00;
                15'h5558: d <= 8'h45; 15'h5559: d <= 8'h35; 15'h555A: d <= 8'hAA; 15'h555B: d <= 8'h00;
                15'h555C: d <= 8'h00; 15'h555D: d <= 8'h00; 15'h555E: d <= 8'h00; 15'h555F: d <= 8'h00;
                15'h5560: d <= 8'h00; 15'h5561: d <= 8'h00; 15'h5562: d <= 8'h00; 15'h5563: d <= 8'h00;
                15'h5564: d <= 8'h00; 15'h5565: d <= 8'h00; 15'h5566: d <= 8'h00; 15'h5567: d <= 8'h00;
                15'h5568: d <= 8'h00; 15'h5569: d <= 8'h00; 15'h556A: d <= 8'h00; 15'h556B: d <= 8'h00;
                15'h556C: d <= 8'h00; 15'h556D: d <= 8'h00; 15'h556E: d <= 8'h00; 15'h556F: d <= 8'h00;
                15'h5570: d <= 8'h00; 15'h5571: d <= 8'h00; 15'h5572: d <= 8'h00; 15'h5573: d <= 8'h00;
                15'h5574: d <= 8'h00; 15'h5575: d <= 8'h00; 15'h5576: d <= 8'h00; 15'h5577: d <= 8'h00;
                15'h5578: d <= 8'h00; 15'h5579: d <= 8'h00; 15'h557A: d <= 8'h00; 15'h557B: d <= 8'h00;
                15'h557C: d <= 8'h00; 15'h557D: d <= 8'h00; 15'h557E: d <= 8'h00; 15'h557F: d <= 8'hE0;
                15'h5580: d <= 8'h10; 15'h5581: d <= 8'h15; 15'h5582: d <= 8'h1A; 15'h5583: d <= 8'h1F;
                15'h5584: d <= 8'h20; 15'h5585: d <= 8'h25; 15'h5586: d <= 8'h2A; 15'h5587: d <= 8'h2F;
                15'h5588: d <= 8'h34; 15'h5589: d <= 8'h38; 15'h558A: d <= 8'h3C; 15'h558B: d <= 8'h31;
                15'h558C: d <= 8'h39; 15'h558D: d <= 8'h3D; 15'h558E: d <= 8'h32; 15'h558F: d <= 8'h36;
                15'h5590: d <= 8'h3E; 15'h5591: d <= 8'h33; 15'h5592: d <= 8'h37; 15'h5593: d <= 8'h3B;
                15'h5594: d <= 8'h44; 15'h5595: d <= 8'h48; 15'h5596: d <= 8'h4C; 15'h5597: d <= 8'h41;
                15'h5598: d <= 8'h49; 15'h5599: d <= 8'h4D; 15'h559A: d <= 8'h42; 15'h559B: d <= 8'h46;
                15'h559C: d <= 8'h4E; 15'h559D: d <= 8'h43; 15'h559E: d <= 8'h47; 15'h559F: d <= 8'h4B;
                15'h55A0: d <= 8'h50; 15'h55A1: d <= 8'h55; 15'h55A2: d <= 8'h5A; 15'h55A3: d <= 8'h5F;
                15'h55A4: d <= 8'h60; 15'h55A5: d <= 8'h65; 15'h55A6: d <= 8'h6A; 15'h55A7: d <= 8'h6F;
                15'h55A8: d <= 8'h74; 15'h55A9: d <= 8'h78; 15'h55AA: d <= 8'h7C; 15'h55AB: d <= 8'h71;
                15'h55AC: d <= 8'h79; 15'h55AD: d <= 8'h7D; 15'h55AE: d <= 8'h72; 15'h55AF: d <= 8'h76;
                15'h55B0: d <= 8'h7E; 15'h55B1: d <= 8'h73; 15'h55B2: d <= 8'h77; 15'h55B3: d <= 8'h7B;
                15'h55B4: d <= 8'h84; 15'h55B5: d <= 8'h88; 15'h55B6: d <= 8'h8C; 15'h55B7: d <= 8'h81;
                15'h55B8: d <= 8'h89; 15'h55B9: d <= 8'h8D; 15'h55BA: d <= 8'h82; 15'h55BB: d <= 8'h86;
                15'h55BC: d <= 8'h8E; 15'h55BD: d <= 8'h83; 15'h55BE: d <= 8'h87; 15'h55BF: d <= 8'h8B;
                15'h55C0: d <= 8'h90; 15'h55C1: d <= 8'h95; 15'h55C2: d <= 8'h9A; 15'h55C3: d <= 8'h9F;
                15'h55C4: d <= 8'hA4; 15'h55C5: d <= 8'hA8; 15'h55C6: d <= 8'hAC; 15'h55C7: d <= 8'hA1;
                15'h55C8: d <= 8'hA9; 15'h55C9: d <= 8'hAD; 15'h55CA: d <= 8'hA2; 15'h55CB: d <= 8'hA6;
                15'h55CC: d <= 8'hAE; 15'h55CD: d <= 8'hA3; 15'h55CE: d <= 8'hA7; 15'h55CF: d <= 8'hAB;
                15'h55D0: d <= 8'hB4; 15'h55D1: d <= 8'hB8; 15'h55D2: d <= 8'hBC; 15'h55D3: d <= 8'hB1;
                15'h55D4: d <= 8'hB9; 15'h55D5: d <= 8'hBD; 15'h55D6: d <= 8'hB2; 15'h55D7: d <= 8'hB6;
                15'h55D8: d <= 8'hBE; 15'h55D9: d <= 8'hB3; 15'h55DA: d <= 8'hB7; 15'h55DB: d <= 8'hBB;
                15'h55DC: d <= 8'hC4; 15'h55DD: d <= 8'hC8; 15'h55DE: d <= 8'hCC; 15'h55DF: d <= 8'hC1;
                15'h55E0: d <= 8'hC9; 15'h55E1: d <= 8'hCD; 15'h55E2: d <= 8'hC2; 15'h55E3: d <= 8'hC6;
                15'h55E4: d <= 8'hCE; 15'h55E5: d <= 8'hC3; 15'h55E6: d <= 8'hC7; 15'h55E7: d <= 8'hCB;
                15'h55E8: d <= 8'hC0; 15'h55E9: d <= 8'hC5; 15'h55EA: d <= 8'hCA; 15'h55EB: d <= 8'hCF;
                15'h55EC: d <= 8'hD0; 15'h55ED: d <= 8'hD5; 15'h55EE: d <= 8'hDA; 15'h55EF: d <= 8'hDF;
                15'h55F0: d <= 8'h74; 15'h55F1: d <= 8'h78; 15'h55F2: d <= 8'h7C; 15'h55F3: d <= 8'h71;
                15'h55F4: d <= 8'h79; 15'h55F5: d <= 8'h7D; 15'h55F6: d <= 8'h72; 15'h55F7: d <= 8'h76;
                15'h55F8: d <= 8'h7E; 15'h55F9: d <= 8'h73; 15'h55FA: d <= 8'h77; 15'h55FB: d <= 8'h7B;
                15'h55FC: d <= 8'hA0; 15'h55FD: d <= 8'hA5; 15'h55FE: d <= 8'hAA; 15'h55FF: d <= 8'hAF;
                15'h5600: d <= 8'h00; 15'h5601: d <= 8'h00; 15'h5602: d <= 8'h00; 15'h5603: d <= 8'h00;
                15'h5604: d <= 8'h00; 15'h5605: d <= 8'h00; 15'h5606: d <= 8'h00; 15'h5607: d <= 8'h00;
                15'h5608: d <= 8'h00; 15'h5609: d <= 8'h00; 15'h560A: d <= 8'h00; 15'h560B: d <= 8'h00;
                15'h560C: d <= 8'h00; 15'h560D: d <= 8'h00; 15'h560E: d <= 8'h00; 15'h560F: d <= 8'h00;
                15'h5610: d <= 8'h00; 15'h5611: d <= 8'h00; 15'h5612: d <= 8'h00; 15'h5613: d <= 8'h00;
                15'h5614: d <= 8'h00; 15'h5615: d <= 8'h00; 15'h5616: d <= 8'h00; 15'h5617: d <= 8'h00;
                15'h5618: d <= 8'h00; 15'h5619: d <= 8'h00; 15'h561A: d <= 8'h00; 15'h561B: d <= 8'h00;
                15'h561C: d <= 8'h00; 15'h561D: d <= 8'h00; 15'h561E: d <= 8'h00; 15'h561F: d <= 8'h00;
                15'h5620: d <= 8'h00; 15'h5621: d <= 8'h00; 15'h5622: d <= 8'h00; 15'h5623: d <= 8'h00;
                15'h5624: d <= 8'h00; 15'h5625: d <= 8'h00; 15'h5626: d <= 8'h00; 15'h5627: d <= 8'h00;
                15'h5628: d <= 8'h00; 15'h5629: d <= 8'h00; 15'h562A: d <= 8'h00; 15'h562B: d <= 8'h00;
                15'h562C: d <= 8'h00; 15'h562D: d <= 8'h00; 15'h562E: d <= 8'h00; 15'h562F: d <= 8'hAF;
                15'h5630: d <= 8'h00; 15'h5631: d <= 8'h00; 15'h5632: d <= 8'h00; 15'h5633: d <= 8'h00;
                15'h5634: d <= 8'h00; 15'h5635: d <= 8'h00; 15'h5636: d <= 8'h00; 15'h5637: d <= 8'h00;
                15'h5638: d <= 8'h00; 15'h5639: d <= 8'h00; 15'h563A: d <= 8'h00; 15'h563B: d <= 8'h00;
                15'h563C: d <= 8'h00; 15'h563D: d <= 8'h00; 15'h563E: d <= 8'h00; 15'h563F: d <= 8'h00;
                15'h5640: d <= 8'h00; 15'h5641: d <= 8'h00; 15'h5642: d <= 8'h00; 15'h5643: d <= 8'h00;
                15'h5644: d <= 8'h00; 15'h5645: d <= 8'h00; 15'h5646: d <= 8'h00; 15'h5647: d <= 8'h00;
                15'h5648: d <= 8'h00; 15'h5649: d <= 8'h00; 15'h564A: d <= 8'h00; 15'h564B: d <= 8'h00;
                15'h564C: d <= 8'h00; 15'h564D: d <= 8'h00; 15'h564E: d <= 8'h00; 15'h564F: d <= 8'h00;
                15'h5650: d <= 8'h00; 15'h5651: d <= 8'h00; 15'h5652: d <= 8'h00; 15'h5653: d <= 8'h00;
                15'h5654: d <= 8'h00; 15'h5655: d <= 8'h00; 15'h5656: d <= 8'h00; 15'h5657: d <= 8'h00;
                15'h5658: d <= 8'h45; 15'h5659: d <= 8'h35; 15'h565A: d <= 8'hAA; 15'h565B: d <= 8'h00;
                15'h565C: d <= 8'h00; 15'h565D: d <= 8'h00; 15'h565E: d <= 8'h00; 15'h565F: d <= 8'h00;
                15'h5660: d <= 8'h00; 15'h5661: d <= 8'h00; 15'h5662: d <= 8'h00; 15'h5663: d <= 8'h00;
                15'h5664: d <= 8'h00; 15'h5665: d <= 8'h00; 15'h5666: d <= 8'h00; 15'h5667: d <= 8'h00;
                15'h5668: d <= 8'h00; 15'h5669: d <= 8'h00; 15'h566A: d <= 8'h00; 15'h566B: d <= 8'h00;
                15'h566C: d <= 8'h00; 15'h566D: d <= 8'h00; 15'h566E: d <= 8'h00; 15'h566F: d <= 8'h00;
                15'h5670: d <= 8'h00; 15'h5671: d <= 8'h00; 15'h5672: d <= 8'h00; 15'h5673: d <= 8'h00;
                15'h5674: d <= 8'h00; 15'h5675: d <= 8'h00; 15'h5676: d <= 8'h00; 15'h5677: d <= 8'h00;
                15'h5678: d <= 8'h00; 15'h5679: d <= 8'h00; 15'h567A: d <= 8'h00; 15'h567B: d <= 8'h00;
                15'h567C: d <= 8'h00; 15'h567D: d <= 8'h00; 15'h567E: d <= 8'h00; 15'h567F: d <= 8'hE0;
                15'h5680: d <= 8'h10; 15'h5681: d <= 8'h15; 15'h5682: d <= 8'h1A; 15'h5683: d <= 8'h1F;
                15'h5684: d <= 8'h20; 15'h5685: d <= 8'h25; 15'h5686: d <= 8'h2A; 15'h5687: d <= 8'h2F;
                15'h5688: d <= 8'h34; 15'h5689: d <= 8'h38; 15'h568A: d <= 8'h3C; 15'h568B: d <= 8'h31;
                15'h568C: d <= 8'h39; 15'h568D: d <= 8'h3D; 15'h568E: d <= 8'h32; 15'h568F: d <= 8'h36;
                15'h5690: d <= 8'h3E; 15'h5691: d <= 8'h33; 15'h5692: d <= 8'h37; 15'h5693: d <= 8'h3B;
                15'h5694: d <= 8'h44; 15'h5695: d <= 8'h48; 15'h5696: d <= 8'h4C; 15'h5697: d <= 8'h41;
                15'h5698: d <= 8'h49; 15'h5699: d <= 8'h4D; 15'h569A: d <= 8'h42; 15'h569B: d <= 8'h46;
                15'h569C: d <= 8'h4E; 15'h569D: d <= 8'h43; 15'h569E: d <= 8'h47; 15'h569F: d <= 8'h4B;
                15'h56A0: d <= 8'h50; 15'h56A1: d <= 8'h55; 15'h56A2: d <= 8'h5A; 15'h56A3: d <= 8'h5F;
                15'h56A4: d <= 8'h60; 15'h56A5: d <= 8'h65; 15'h56A6: d <= 8'h6A; 15'h56A7: d <= 8'h6F;
                15'h56A8: d <= 8'h74; 15'h56A9: d <= 8'h78; 15'h56AA: d <= 8'h7C; 15'h56AB: d <= 8'h71;
                15'h56AC: d <= 8'h79; 15'h56AD: d <= 8'h7D; 15'h56AE: d <= 8'h72; 15'h56AF: d <= 8'h76;
                15'h56B0: d <= 8'h7E; 15'h56B1: d <= 8'h73; 15'h56B2: d <= 8'h77; 15'h56B3: d <= 8'h7B;
                15'h56B4: d <= 8'h84; 15'h56B5: d <= 8'h88; 15'h56B6: d <= 8'h8C; 15'h56B7: d <= 8'h81;
                15'h56B8: d <= 8'h89; 15'h56B9: d <= 8'h8D; 15'h56BA: d <= 8'h82; 15'h56BB: d <= 8'h86;
                15'h56BC: d <= 8'h8E; 15'h56BD: d <= 8'h83; 15'h56BE: d <= 8'h87; 15'h56BF: d <= 8'h8B;
                15'h56C0: d <= 8'h90; 15'h56C1: d <= 8'h95; 15'h56C2: d <= 8'h9A; 15'h56C3: d <= 8'h9F;
                15'h56C4: d <= 8'hA4; 15'h56C5: d <= 8'hA8; 15'h56C6: d <= 8'hAC; 15'h56C7: d <= 8'hA1;
                15'h56C8: d <= 8'hA9; 15'h56C9: d <= 8'hAD; 15'h56CA: d <= 8'hA2; 15'h56CB: d <= 8'hA6;
                15'h56CC: d <= 8'hAE; 15'h56CD: d <= 8'hA3; 15'h56CE: d <= 8'hA7; 15'h56CF: d <= 8'hAB;
                15'h56D0: d <= 8'hB4; 15'h56D1: d <= 8'hB8; 15'h56D2: d <= 8'hBC; 15'h56D3: d <= 8'hB1;
                15'h56D4: d <= 8'hB9; 15'h56D5: d <= 8'hBD; 15'h56D6: d <= 8'hB2; 15'h56D7: d <= 8'hB6;
                15'h56D8: d <= 8'hBE; 15'h56D9: d <= 8'hB3; 15'h56DA: d <= 8'hB7; 15'h56DB: d <= 8'hBB;
                15'h56DC: d <= 8'hC4; 15'h56DD: d <= 8'hC8; 15'h56DE: d <= 8'hCC; 15'h56DF: d <= 8'hC1;
                15'h56E0: d <= 8'hC9; 15'h56E1: d <= 8'hCD; 15'h56E2: d <= 8'hC2; 15'h56E3: d <= 8'hC6;
                15'h56E4: d <= 8'hCE; 15'h56E5: d <= 8'hC3; 15'h56E6: d <= 8'hC7; 15'h56E7: d <= 8'hCB;
                15'h56E8: d <= 8'hC0; 15'h56E9: d <= 8'hC5; 15'h56EA: d <= 8'hCA; 15'h56EB: d <= 8'hCF;
                15'h56EC: d <= 8'hD0; 15'h56ED: d <= 8'hD5; 15'h56EE: d <= 8'hDA; 15'h56EF: d <= 8'hDF;
                15'h56F0: d <= 8'h74; 15'h56F1: d <= 8'h78; 15'h56F2: d <= 8'h7C; 15'h56F3: d <= 8'h71;
                15'h56F4: d <= 8'h79; 15'h56F5: d <= 8'h7D; 15'h56F6: d <= 8'h72; 15'h56F7: d <= 8'h76;
                15'h56F8: d <= 8'h7E; 15'h56F9: d <= 8'h73; 15'h56FA: d <= 8'h77; 15'h56FB: d <= 8'h7B;
                15'h56FC: d <= 8'hA0; 15'h56FD: d <= 8'hA5; 15'h56FE: d <= 8'hAA; 15'h56FF: d <= 8'hAF;
                15'h5700: d <= 8'h00; 15'h5701: d <= 8'h00; 15'h5702: d <= 8'h00; 15'h5703: d <= 8'h00;
                15'h5704: d <= 8'h00; 15'h5705: d <= 8'h00; 15'h5706: d <= 8'h00; 15'h5707: d <= 8'h00;
                15'h5708: d <= 8'h00; 15'h5709: d <= 8'h00; 15'h570A: d <= 8'h00; 15'h570B: d <= 8'h00;
                15'h570C: d <= 8'h00; 15'h570D: d <= 8'h00; 15'h570E: d <= 8'h00; 15'h570F: d <= 8'h00;
                15'h5710: d <= 8'h00; 15'h5711: d <= 8'h00; 15'h5712: d <= 8'h00; 15'h5713: d <= 8'h00;
                15'h5714: d <= 8'h00; 15'h5715: d <= 8'h00; 15'h5716: d <= 8'h00; 15'h5717: d <= 8'h00;
                15'h5718: d <= 8'h00; 15'h5719: d <= 8'h00; 15'h571A: d <= 8'h00; 15'h571B: d <= 8'h00;
                15'h571C: d <= 8'h00; 15'h571D: d <= 8'h00; 15'h571E: d <= 8'h00; 15'h571F: d <= 8'h00;
                15'h5720: d <= 8'h00; 15'h5721: d <= 8'h00; 15'h5722: d <= 8'h00; 15'h5723: d <= 8'h00;
                15'h5724: d <= 8'h00; 15'h5725: d <= 8'h00; 15'h5726: d <= 8'h00; 15'h5727: d <= 8'h00;
                15'h5728: d <= 8'h00; 15'h5729: d <= 8'h00; 15'h572A: d <= 8'h00; 15'h572B: d <= 8'h00;
                15'h572C: d <= 8'h00; 15'h572D: d <= 8'h00; 15'h572E: d <= 8'h00; 15'h572F: d <= 8'hAF;
                15'h5730: d <= 8'h00; 15'h5731: d <= 8'h00; 15'h5732: d <= 8'h00; 15'h5733: d <= 8'h00;
                15'h5734: d <= 8'h00; 15'h5735: d <= 8'h00; 15'h5736: d <= 8'h00; 15'h5737: d <= 8'h00;
                15'h5738: d <= 8'h00; 15'h5739: d <= 8'h00; 15'h573A: d <= 8'h00; 15'h573B: d <= 8'h00;
                15'h573C: d <= 8'h00; 15'h573D: d <= 8'h00; 15'h573E: d <= 8'h00; 15'h573F: d <= 8'h00;
                15'h5740: d <= 8'h00; 15'h5741: d <= 8'h00; 15'h5742: d <= 8'h00; 15'h5743: d <= 8'h00;
                15'h5744: d <= 8'h00; 15'h5745: d <= 8'h00; 15'h5746: d <= 8'h00; 15'h5747: d <= 8'h00;
                15'h5748: d <= 8'h00; 15'h5749: d <= 8'h00; 15'h574A: d <= 8'h00; 15'h574B: d <= 8'h00;
                15'h574C: d <= 8'h00; 15'h574D: d <= 8'h00; 15'h574E: d <= 8'h00; 15'h574F: d <= 8'h00;
                15'h5750: d <= 8'h00; 15'h5751: d <= 8'h00; 15'h5752: d <= 8'h00; 15'h5753: d <= 8'h00;
                15'h5754: d <= 8'h00; 15'h5755: d <= 8'h00; 15'h5756: d <= 8'h00; 15'h5757: d <= 8'h00;
                15'h5758: d <= 8'h45; 15'h5759: d <= 8'h35; 15'h575A: d <= 8'hAA; 15'h575B: d <= 8'h00;
                15'h575C: d <= 8'h00; 15'h575D: d <= 8'h00; 15'h575E: d <= 8'h00; 15'h575F: d <= 8'h00;
                15'h5760: d <= 8'h00; 15'h5761: d <= 8'h00; 15'h5762: d <= 8'h00; 15'h5763: d <= 8'h00;
                15'h5764: d <= 8'h00; 15'h5765: d <= 8'h00; 15'h5766: d <= 8'h00; 15'h5767: d <= 8'h00;
                15'h5768: d <= 8'h00; 15'h5769: d <= 8'h00; 15'h576A: d <= 8'h00; 15'h576B: d <= 8'h00;
                15'h576C: d <= 8'h00; 15'h576D: d <= 8'h00; 15'h576E: d <= 8'h00; 15'h576F: d <= 8'h00;
                15'h5770: d <= 8'h00; 15'h5771: d <= 8'h00; 15'h5772: d <= 8'h00; 15'h5773: d <= 8'h00;
                15'h5774: d <= 8'h00; 15'h5775: d <= 8'h00; 15'h5776: d <= 8'h00; 15'h5777: d <= 8'h00;
                15'h5778: d <= 8'h00; 15'h5779: d <= 8'h00; 15'h577A: d <= 8'h00; 15'h577B: d <= 8'h00;
                15'h577C: d <= 8'h00; 15'h577D: d <= 8'h00; 15'h577E: d <= 8'h00; 15'h577F: d <= 8'hE0;
                15'h5780: d <= 8'h10; 15'h5781: d <= 8'h15; 15'h5782: d <= 8'h1A; 15'h5783: d <= 8'h1F;
                15'h5784: d <= 8'h20; 15'h5785: d <= 8'h25; 15'h5786: d <= 8'h2A; 15'h5787: d <= 8'h2F;
                15'h5788: d <= 8'h34; 15'h5789: d <= 8'h38; 15'h578A: d <= 8'h3C; 15'h578B: d <= 8'h31;
                15'h578C: d <= 8'h39; 15'h578D: d <= 8'h3D; 15'h578E: d <= 8'h32; 15'h578F: d <= 8'h36;
                15'h5790: d <= 8'h3E; 15'h5791: d <= 8'h33; 15'h5792: d <= 8'h37; 15'h5793: d <= 8'h3B;
                15'h5794: d <= 8'h44; 15'h5795: d <= 8'h48; 15'h5796: d <= 8'h4C; 15'h5797: d <= 8'h41;
                15'h5798: d <= 8'h49; 15'h5799: d <= 8'h4D; 15'h579A: d <= 8'h42; 15'h579B: d <= 8'h46;
                15'h579C: d <= 8'h4E; 15'h579D: d <= 8'h43; 15'h579E: d <= 8'h47; 15'h579F: d <= 8'h4B;
                15'h57A0: d <= 8'h50; 15'h57A1: d <= 8'h55; 15'h57A2: d <= 8'h5A; 15'h57A3: d <= 8'h5F;
                15'h57A4: d <= 8'h60; 15'h57A5: d <= 8'h65; 15'h57A6: d <= 8'h6A; 15'h57A7: d <= 8'h6F;
                15'h57A8: d <= 8'h74; 15'h57A9: d <= 8'h78; 15'h57AA: d <= 8'h7C; 15'h57AB: d <= 8'h71;
                15'h57AC: d <= 8'h79; 15'h57AD: d <= 8'h7D; 15'h57AE: d <= 8'h72; 15'h57AF: d <= 8'h76;
                15'h57B0: d <= 8'h7E; 15'h57B1: d <= 8'h73; 15'h57B2: d <= 8'h77; 15'h57B3: d <= 8'h7B;
                15'h57B4: d <= 8'h84; 15'h57B5: d <= 8'h88; 15'h57B6: d <= 8'h8C; 15'h57B7: d <= 8'h81;
                15'h57B8: d <= 8'h89; 15'h57B9: d <= 8'h8D; 15'h57BA: d <= 8'h82; 15'h57BB: d <= 8'h86;
                15'h57BC: d <= 8'h8E; 15'h57BD: d <= 8'h83; 15'h57BE: d <= 8'h87; 15'h57BF: d <= 8'h8B;
                15'h57C0: d <= 8'h90; 15'h57C1: d <= 8'h95; 15'h57C2: d <= 8'h9A; 15'h57C3: d <= 8'h9F;
                15'h57C4: d <= 8'hA4; 15'h57C5: d <= 8'hA8; 15'h57C6: d <= 8'hAC; 15'h57C7: d <= 8'hA1;
                15'h57C8: d <= 8'hA9; 15'h57C9: d <= 8'hAD; 15'h57CA: d <= 8'hA2; 15'h57CB: d <= 8'hA6;
                15'h57CC: d <= 8'hAE; 15'h57CD: d <= 8'hA3; 15'h57CE: d <= 8'hA7; 15'h57CF: d <= 8'hAB;
                15'h57D0: d <= 8'hB4; 15'h57D1: d <= 8'hB8; 15'h57D2: d <= 8'hBC; 15'h57D3: d <= 8'hB1;
                15'h57D4: d <= 8'hB9; 15'h57D5: d <= 8'hBD; 15'h57D6: d <= 8'hB2; 15'h57D7: d <= 8'hB6;
                15'h57D8: d <= 8'hBE; 15'h57D9: d <= 8'hB3; 15'h57DA: d <= 8'hB7; 15'h57DB: d <= 8'hBB;
                15'h57DC: d <= 8'hC4; 15'h57DD: d <= 8'hC8; 15'h57DE: d <= 8'hCC; 15'h57DF: d <= 8'hC1;
                15'h57E0: d <= 8'hC9; 15'h57E1: d <= 8'hCD; 15'h57E2: d <= 8'hC2; 15'h57E3: d <= 8'hC6;
                15'h57E4: d <= 8'hCE; 15'h57E5: d <= 8'hC3; 15'h57E6: d <= 8'hC7; 15'h57E7: d <= 8'hCB;
                15'h57E8: d <= 8'hC0; 15'h57E9: d <= 8'hC5; 15'h57EA: d <= 8'hCA; 15'h57EB: d <= 8'hCF;
                15'h57EC: d <= 8'hD0; 15'h57ED: d <= 8'hD5; 15'h57EE: d <= 8'hDA; 15'h57EF: d <= 8'hDF;
                15'h57F0: d <= 8'h74; 15'h57F1: d <= 8'h78; 15'h57F2: d <= 8'h7C; 15'h57F3: d <= 8'h71;
                15'h57F4: d <= 8'h79; 15'h57F5: d <= 8'h7D; 15'h57F6: d <= 8'h72; 15'h57F7: d <= 8'h76;
                15'h57F8: d <= 8'h7E; 15'h57F9: d <= 8'h73; 15'h57FA: d <= 8'h77; 15'h57FB: d <= 8'h7B;
                15'h57FC: d <= 8'hA0; 15'h57FD: d <= 8'hA5; 15'h57FE: d <= 8'hAA; 15'h57FF: d <= 8'hAF;
                15'h5800: d <= 8'h00; 15'h5801: d <= 8'h00; 15'h5802: d <= 8'h00; 15'h5803: d <= 8'h00;
                15'h5804: d <= 8'h00; 15'h5805: d <= 8'h00; 15'h5806: d <= 8'h00; 15'h5807: d <= 8'h00;
                15'h5808: d <= 8'h00; 15'h5809: d <= 8'h00; 15'h580A: d <= 8'h00; 15'h580B: d <= 8'h00;
                15'h580C: d <= 8'h00; 15'h580D: d <= 8'h00; 15'h580E: d <= 8'h00; 15'h580F: d <= 8'h00;
                15'h5810: d <= 8'h00; 15'h5811: d <= 8'h00; 15'h5812: d <= 8'h00; 15'h5813: d <= 8'h00;
                15'h5814: d <= 8'h00; 15'h5815: d <= 8'h00; 15'h5816: d <= 8'h00; 15'h5817: d <= 8'h00;
                15'h5818: d <= 8'h00; 15'h5819: d <= 8'h00; 15'h581A: d <= 8'h00; 15'h581B: d <= 8'h00;
                15'h581C: d <= 8'h00; 15'h581D: d <= 8'h00; 15'h581E: d <= 8'h00; 15'h581F: d <= 8'h00;
                15'h5820: d <= 8'h00; 15'h5821: d <= 8'h00; 15'h5822: d <= 8'h00; 15'h5823: d <= 8'h00;
                15'h5824: d <= 8'h00; 15'h5825: d <= 8'h00; 15'h5826: d <= 8'h00; 15'h5827: d <= 8'h00;
                15'h5828: d <= 8'h00; 15'h5829: d <= 8'h00; 15'h582A: d <= 8'h00; 15'h582B: d <= 8'h00;
                15'h582C: d <= 8'h00; 15'h582D: d <= 8'h00; 15'h582E: d <= 8'h00; 15'h582F: d <= 8'h7B;
                15'h5830: d <= 8'h00; 15'h5831: d <= 8'h00; 15'h5832: d <= 8'h00; 15'h5833: d <= 8'h00;
                15'h5834: d <= 8'h00; 15'h5835: d <= 8'h00; 15'h5836: d <= 8'h00; 15'h5837: d <= 8'h00;
                15'h5838: d <= 8'h00; 15'h5839: d <= 8'h00; 15'h583A: d <= 8'h00; 15'h583B: d <= 8'h00;
                15'h583C: d <= 8'h00; 15'h583D: d <= 8'h00; 15'h583E: d <= 8'h00; 15'h583F: d <= 8'h00;
                15'h5840: d <= 8'h00; 15'h5841: d <= 8'h00; 15'h5842: d <= 8'h00; 15'h5843: d <= 8'h00;
                15'h5844: d <= 8'h00; 15'h5845: d <= 8'h00; 15'h5846: d <= 8'h00; 15'h5847: d <= 8'h00;
                15'h5848: d <= 8'h00; 15'h5849: d <= 8'h00; 15'h584A: d <= 8'h00; 15'h584B: d <= 8'h00;
                15'h584C: d <= 8'h00; 15'h584D: d <= 8'h00; 15'h584E: d <= 8'h00; 15'h584F: d <= 8'h00;
                15'h5850: d <= 8'h00; 15'h5851: d <= 8'h00; 15'h5852: d <= 8'h00; 15'h5853: d <= 8'h00;
                15'h5854: d <= 8'h00; 15'h5855: d <= 8'h00; 15'h5856: d <= 8'h00; 15'h5857: d <= 8'h00;
                15'h5858: d <= 8'h45; 15'h5859: d <= 8'h35; 15'h585A: d <= 8'h32; 15'h585B: d <= 8'h00;
                15'h585C: d <= 8'h00; 15'h585D: d <= 8'h00; 15'h585E: d <= 8'h00; 15'h585F: d <= 8'h00;
                15'h5860: d <= 8'h00; 15'h5861: d <= 8'h00; 15'h5862: d <= 8'h00; 15'h5863: d <= 8'h00;
                15'h5864: d <= 8'h00; 15'h5865: d <= 8'h00; 15'h5866: d <= 8'h00; 15'h5867: d <= 8'h00;
                15'h5868: d <= 8'h00; 15'h5869: d <= 8'h00; 15'h586A: d <= 8'h00; 15'h586B: d <= 8'h00;
                15'h586C: d <= 8'h00; 15'h586D: d <= 8'h00; 15'h586E: d <= 8'h00; 15'h586F: d <= 8'h00;
                15'h5870: d <= 8'h00; 15'h5871: d <= 8'h00; 15'h5872: d <= 8'h00; 15'h5873: d <= 8'h00;
                15'h5874: d <= 8'h00; 15'h5875: d <= 8'h00; 15'h5876: d <= 8'h00; 15'h5877: d <= 8'h00;
                15'h5878: d <= 8'h00; 15'h5879: d <= 8'h00; 15'h587A: d <= 8'h00; 15'h587B: d <= 8'h00;
                15'h587C: d <= 8'h00; 15'h587D: d <= 8'h00; 15'h587E: d <= 8'h00; 15'h587F: d <= 8'hE0;
                15'h5880: d <= 8'h10; 15'h5881: d <= 8'h15; 15'h5882: d <= 8'h1A; 15'h5883: d <= 8'h1F;
                15'h5884: d <= 8'h20; 15'h5885: d <= 8'h25; 15'h5886: d <= 8'h2A; 15'h5887: d <= 8'h2F;
                15'h5888: d <= 8'h34; 15'h5889: d <= 8'h38; 15'h588A: d <= 8'h3C; 15'h588B: d <= 8'h31;
                15'h588C: d <= 8'h39; 15'h588D: d <= 8'h3D; 15'h588E: d <= 8'h32; 15'h588F: d <= 8'h36;
                15'h5890: d <= 8'h3E; 15'h5891: d <= 8'h33; 15'h5892: d <= 8'h37; 15'h5893: d <= 8'h3B;
                15'h5894: d <= 8'h44; 15'h5895: d <= 8'h48; 15'h5896: d <= 8'h4C; 15'h5897: d <= 8'h41;
                15'h5898: d <= 8'h49; 15'h5899: d <= 8'h4D; 15'h589A: d <= 8'h42; 15'h589B: d <= 8'h46;
                15'h589C: d <= 8'h4E; 15'h589D: d <= 8'h43; 15'h589E: d <= 8'h47; 15'h589F: d <= 8'h4B;
                15'h58A0: d <= 8'h50; 15'h58A1: d <= 8'h55; 15'h58A2: d <= 8'h5A; 15'h58A3: d <= 8'h5F;
                15'h58A4: d <= 8'h60; 15'h58A5: d <= 8'h65; 15'h58A6: d <= 8'h6A; 15'h58A7: d <= 8'h6F;
                15'h58A8: d <= 8'h74; 15'h58A9: d <= 8'h78; 15'h58AA: d <= 8'h7C; 15'h58AB: d <= 8'h71;
                15'h58AC: d <= 8'h79; 15'h58AD: d <= 8'h7D; 15'h58AE: d <= 8'h72; 15'h58AF: d <= 8'h76;
                15'h58B0: d <= 8'h7E; 15'h58B1: d <= 8'h73; 15'h58B2: d <= 8'h77; 15'h58B3: d <= 8'h7B;
                15'h58B4: d <= 8'h84; 15'h58B5: d <= 8'h88; 15'h58B6: d <= 8'h8C; 15'h58B7: d <= 8'h81;
                15'h58B8: d <= 8'h89; 15'h58B9: d <= 8'h8D; 15'h58BA: d <= 8'h82; 15'h58BB: d <= 8'h86;
                15'h58BC: d <= 8'h8E; 15'h58BD: d <= 8'h83; 15'h58BE: d <= 8'h87; 15'h58BF: d <= 8'h8B;
                15'h58C0: d <= 8'h90; 15'h58C1: d <= 8'h95; 15'h58C2: d <= 8'h9A; 15'h58C3: d <= 8'h9F;
                15'h58C4: d <= 8'hA4; 15'h58C5: d <= 8'hA8; 15'h58C6: d <= 8'hAC; 15'h58C7: d <= 8'hA1;
                15'h58C8: d <= 8'hA9; 15'h58C9: d <= 8'hAD; 15'h58CA: d <= 8'hA2; 15'h58CB: d <= 8'hA6;
                15'h58CC: d <= 8'hAE; 15'h58CD: d <= 8'hA3; 15'h58CE: d <= 8'hA7; 15'h58CF: d <= 8'hAB;
                15'h58D0: d <= 8'hB4; 15'h58D1: d <= 8'hB8; 15'h58D2: d <= 8'hBC; 15'h58D3: d <= 8'hB1;
                15'h58D4: d <= 8'hB9; 15'h58D5: d <= 8'hBD; 15'h58D6: d <= 8'hB2; 15'h58D7: d <= 8'hB6;
                15'h58D8: d <= 8'hBE; 15'h58D9: d <= 8'hB3; 15'h58DA: d <= 8'hB7; 15'h58DB: d <= 8'hBB;
                15'h58DC: d <= 8'hC4; 15'h58DD: d <= 8'hC8; 15'h58DE: d <= 8'hCC; 15'h58DF: d <= 8'hC1;
                15'h58E0: d <= 8'hC9; 15'h58E1: d <= 8'hCD; 15'h58E2: d <= 8'hC2; 15'h58E3: d <= 8'hC6;
                15'h58E4: d <= 8'hCE; 15'h58E5: d <= 8'hC3; 15'h58E6: d <= 8'hC7; 15'h58E7: d <= 8'hCB;
                15'h58E8: d <= 8'hC0; 15'h58E9: d <= 8'hC5; 15'h58EA: d <= 8'hCA; 15'h58EB: d <= 8'hCF;
                15'h58EC: d <= 8'hD0; 15'h58ED: d <= 8'hD5; 15'h58EE: d <= 8'hDA; 15'h58EF: d <= 8'hDF;
                15'h58F0: d <= 8'h74; 15'h58F1: d <= 8'h78; 15'h58F2: d <= 8'h7C; 15'h58F3: d <= 8'h71;
                15'h58F4: d <= 8'h79; 15'h58F5: d <= 8'h7D; 15'h58F6: d <= 8'h72; 15'h58F7: d <= 8'h76;
                15'h58F8: d <= 8'h7E; 15'h58F9: d <= 8'h73; 15'h58FA: d <= 8'h77; 15'h58FB: d <= 8'h7B;
                15'h58FC: d <= 8'hA0; 15'h58FD: d <= 8'hA5; 15'h58FE: d <= 8'hAA; 15'h58FF: d <= 8'hAF;
                15'h5900: d <= 8'h00; 15'h5901: d <= 8'h00; 15'h5902: d <= 8'h00; 15'h5903: d <= 8'h00;
                15'h5904: d <= 8'h00; 15'h5905: d <= 8'h00; 15'h5906: d <= 8'h00; 15'h5907: d <= 8'h00;
                15'h5908: d <= 8'h00; 15'h5909: d <= 8'h00; 15'h590A: d <= 8'h00; 15'h590B: d <= 8'h00;
                15'h590C: d <= 8'h00; 15'h590D: d <= 8'h00; 15'h590E: d <= 8'h00; 15'h590F: d <= 8'h00;
                15'h5910: d <= 8'h00; 15'h5911: d <= 8'h00; 15'h5912: d <= 8'h00; 15'h5913: d <= 8'h00;
                15'h5914: d <= 8'h00; 15'h5915: d <= 8'h00; 15'h5916: d <= 8'h00; 15'h5917: d <= 8'h00;
                15'h5918: d <= 8'h00; 15'h5919: d <= 8'h00; 15'h591A: d <= 8'h00; 15'h591B: d <= 8'h00;
                15'h591C: d <= 8'h00; 15'h591D: d <= 8'h00; 15'h591E: d <= 8'h00; 15'h591F: d <= 8'h00;
                15'h5920: d <= 8'h00; 15'h5921: d <= 8'h00; 15'h5922: d <= 8'h00; 15'h5923: d <= 8'h00;
                15'h5924: d <= 8'h00; 15'h5925: d <= 8'h00; 15'h5926: d <= 8'h00; 15'h5927: d <= 8'h00;
                15'h5928: d <= 8'h00; 15'h5929: d <= 8'h00; 15'h592A: d <= 8'h00; 15'h592B: d <= 8'h00;
                15'h592C: d <= 8'h00; 15'h592D: d <= 8'h00; 15'h592E: d <= 8'h00; 15'h592F: d <= 8'h7B;
                15'h5930: d <= 8'h00; 15'h5931: d <= 8'h00; 15'h5932: d <= 8'h00; 15'h5933: d <= 8'h00;
                15'h5934: d <= 8'h00; 15'h5935: d <= 8'h00; 15'h5936: d <= 8'h00; 15'h5937: d <= 8'h00;
                15'h5938: d <= 8'h00; 15'h5939: d <= 8'h00; 15'h593A: d <= 8'h00; 15'h593B: d <= 8'h00;
                15'h593C: d <= 8'h00; 15'h593D: d <= 8'h00; 15'h593E: d <= 8'h00; 15'h593F: d <= 8'h00;
                15'h5940: d <= 8'h00; 15'h5941: d <= 8'h00; 15'h5942: d <= 8'h00; 15'h5943: d <= 8'h00;
                15'h5944: d <= 8'h00; 15'h5945: d <= 8'h00; 15'h5946: d <= 8'h00; 15'h5947: d <= 8'h00;
                15'h5948: d <= 8'h00; 15'h5949: d <= 8'h00; 15'h594A: d <= 8'h00; 15'h594B: d <= 8'h00;
                15'h594C: d <= 8'h00; 15'h594D: d <= 8'h00; 15'h594E: d <= 8'h00; 15'h594F: d <= 8'h00;
                15'h5950: d <= 8'h00; 15'h5951: d <= 8'h00; 15'h5952: d <= 8'h00; 15'h5953: d <= 8'h00;
                15'h5954: d <= 8'h00; 15'h5955: d <= 8'h00; 15'h5956: d <= 8'h00; 15'h5957: d <= 8'h00;
                15'h5958: d <= 8'h45; 15'h5959: d <= 8'h35; 15'h595A: d <= 8'h32; 15'h595B: d <= 8'h00;
                15'h595C: d <= 8'h00; 15'h595D: d <= 8'h00; 15'h595E: d <= 8'h00; 15'h595F: d <= 8'h00;
                15'h5960: d <= 8'h00; 15'h5961: d <= 8'h00; 15'h5962: d <= 8'h00; 15'h5963: d <= 8'h00;
                15'h5964: d <= 8'h00; 15'h5965: d <= 8'h00; 15'h5966: d <= 8'h00; 15'h5967: d <= 8'h00;
                15'h5968: d <= 8'h00; 15'h5969: d <= 8'h00; 15'h596A: d <= 8'h00; 15'h596B: d <= 8'h00;
                15'h596C: d <= 8'h00; 15'h596D: d <= 8'h00; 15'h596E: d <= 8'h00; 15'h596F: d <= 8'h00;
                15'h5970: d <= 8'h00; 15'h5971: d <= 8'h00; 15'h5972: d <= 8'h00; 15'h5973: d <= 8'h00;
                15'h5974: d <= 8'h00; 15'h5975: d <= 8'h00; 15'h5976: d <= 8'h00; 15'h5977: d <= 8'h00;
                15'h5978: d <= 8'h00; 15'h5979: d <= 8'h00; 15'h597A: d <= 8'h00; 15'h597B: d <= 8'h00;
                15'h597C: d <= 8'h00; 15'h597D: d <= 8'h00; 15'h597E: d <= 8'h00; 15'h597F: d <= 8'hE0;
                15'h5980: d <= 8'h10; 15'h5981: d <= 8'h15; 15'h5982: d <= 8'h1A; 15'h5983: d <= 8'h1F;
                15'h5984: d <= 8'h20; 15'h5985: d <= 8'h25; 15'h5986: d <= 8'h2A; 15'h5987: d <= 8'h2F;
                15'h5988: d <= 8'h34; 15'h5989: d <= 8'h38; 15'h598A: d <= 8'h3C; 15'h598B: d <= 8'h31;
                15'h598C: d <= 8'h39; 15'h598D: d <= 8'h3D; 15'h598E: d <= 8'h32; 15'h598F: d <= 8'h36;
                15'h5990: d <= 8'h3E; 15'h5991: d <= 8'h33; 15'h5992: d <= 8'h37; 15'h5993: d <= 8'h3B;
                15'h5994: d <= 8'h44; 15'h5995: d <= 8'h48; 15'h5996: d <= 8'h4C; 15'h5997: d <= 8'h41;
                15'h5998: d <= 8'h49; 15'h5999: d <= 8'h4D; 15'h599A: d <= 8'h42; 15'h599B: d <= 8'h46;
                15'h599C: d <= 8'h4E; 15'h599D: d <= 8'h43; 15'h599E: d <= 8'h47; 15'h599F: d <= 8'h4B;
                15'h59A0: d <= 8'h50; 15'h59A1: d <= 8'h55; 15'h59A2: d <= 8'h5A; 15'h59A3: d <= 8'h5F;
                15'h59A4: d <= 8'h60; 15'h59A5: d <= 8'h65; 15'h59A6: d <= 8'h6A; 15'h59A7: d <= 8'h6F;
                15'h59A8: d <= 8'h74; 15'h59A9: d <= 8'h78; 15'h59AA: d <= 8'h7C; 15'h59AB: d <= 8'h71;
                15'h59AC: d <= 8'h79; 15'h59AD: d <= 8'h7D; 15'h59AE: d <= 8'h72; 15'h59AF: d <= 8'h76;
                15'h59B0: d <= 8'h7E; 15'h59B1: d <= 8'h73; 15'h59B2: d <= 8'h77; 15'h59B3: d <= 8'h7B;
                15'h59B4: d <= 8'h84; 15'h59B5: d <= 8'h88; 15'h59B6: d <= 8'h8C; 15'h59B7: d <= 8'h81;
                15'h59B8: d <= 8'h89; 15'h59B9: d <= 8'h8D; 15'h59BA: d <= 8'h82; 15'h59BB: d <= 8'h86;
                15'h59BC: d <= 8'h8E; 15'h59BD: d <= 8'h83; 15'h59BE: d <= 8'h87; 15'h59BF: d <= 8'h8B;
                15'h59C0: d <= 8'h90; 15'h59C1: d <= 8'h95; 15'h59C2: d <= 8'h9A; 15'h59C3: d <= 8'h9F;
                15'h59C4: d <= 8'hA4; 15'h59C5: d <= 8'hA8; 15'h59C6: d <= 8'hAC; 15'h59C7: d <= 8'hA1;
                15'h59C8: d <= 8'hA9; 15'h59C9: d <= 8'hAD; 15'h59CA: d <= 8'hA2; 15'h59CB: d <= 8'hA6;
                15'h59CC: d <= 8'hAE; 15'h59CD: d <= 8'hA3; 15'h59CE: d <= 8'hA7; 15'h59CF: d <= 8'hAB;
                15'h59D0: d <= 8'hB4; 15'h59D1: d <= 8'hB8; 15'h59D2: d <= 8'hBC; 15'h59D3: d <= 8'hB1;
                15'h59D4: d <= 8'hB9; 15'h59D5: d <= 8'hBD; 15'h59D6: d <= 8'hB2; 15'h59D7: d <= 8'hB6;
                15'h59D8: d <= 8'hBE; 15'h59D9: d <= 8'hB3; 15'h59DA: d <= 8'hB7; 15'h59DB: d <= 8'hBB;
                15'h59DC: d <= 8'hC4; 15'h59DD: d <= 8'hC8; 15'h59DE: d <= 8'hCC; 15'h59DF: d <= 8'hC1;
                15'h59E0: d <= 8'hC9; 15'h59E1: d <= 8'hCD; 15'h59E2: d <= 8'hC2; 15'h59E3: d <= 8'hC6;
                15'h59E4: d <= 8'hCE; 15'h59E5: d <= 8'hC3; 15'h59E6: d <= 8'hC7; 15'h59E7: d <= 8'hCB;
                15'h59E8: d <= 8'hC0; 15'h59E9: d <= 8'hC5; 15'h59EA: d <= 8'hCA; 15'h59EB: d <= 8'hCF;
                15'h59EC: d <= 8'hD0; 15'h59ED: d <= 8'hD5; 15'h59EE: d <= 8'hDA; 15'h59EF: d <= 8'hDF;
                15'h59F0: d <= 8'h74; 15'h59F1: d <= 8'h78; 15'h59F2: d <= 8'h7C; 15'h59F3: d <= 8'h71;
                15'h59F4: d <= 8'h79; 15'h59F5: d <= 8'h7D; 15'h59F6: d <= 8'h72; 15'h59F7: d <= 8'h76;
                15'h59F8: d <= 8'h7E; 15'h59F9: d <= 8'h73; 15'h59FA: d <= 8'h77; 15'h59FB: d <= 8'h7B;
                15'h59FC: d <= 8'hA0; 15'h59FD: d <= 8'hA5; 15'h59FE: d <= 8'hAA; 15'h59FF: d <= 8'hAF;
                15'h5A00: d <= 8'h00; 15'h5A01: d <= 8'h00; 15'h5A02: d <= 8'h00; 15'h5A03: d <= 8'h00;
                15'h5A04: d <= 8'h00; 15'h5A05: d <= 8'h00; 15'h5A06: d <= 8'h00; 15'h5A07: d <= 8'h00;
                15'h5A08: d <= 8'h00; 15'h5A09: d <= 8'h00; 15'h5A0A: d <= 8'h00; 15'h5A0B: d <= 8'h00;
                15'h5A0C: d <= 8'h00; 15'h5A0D: d <= 8'h00; 15'h5A0E: d <= 8'h00; 15'h5A0F: d <= 8'h00;
                15'h5A10: d <= 8'h00; 15'h5A11: d <= 8'h00; 15'h5A12: d <= 8'h00; 15'h5A13: d <= 8'h00;
                15'h5A14: d <= 8'h00; 15'h5A15: d <= 8'h00; 15'h5A16: d <= 8'h00; 15'h5A17: d <= 8'h00;
                15'h5A18: d <= 8'h00; 15'h5A19: d <= 8'h00; 15'h5A1A: d <= 8'h00; 15'h5A1B: d <= 8'h00;
                15'h5A1C: d <= 8'h00; 15'h5A1D: d <= 8'h00; 15'h5A1E: d <= 8'h00; 15'h5A1F: d <= 8'h00;
                15'h5A20: d <= 8'h00; 15'h5A21: d <= 8'h00; 15'h5A22: d <= 8'h00; 15'h5A23: d <= 8'h00;
                15'h5A24: d <= 8'h00; 15'h5A25: d <= 8'h00; 15'h5A26: d <= 8'h00; 15'h5A27: d <= 8'h00;
                15'h5A28: d <= 8'h00; 15'h5A29: d <= 8'h00; 15'h5A2A: d <= 8'h00; 15'h5A2B: d <= 8'h00;
                15'h5A2C: d <= 8'h00; 15'h5A2D: d <= 8'h00; 15'h5A2E: d <= 8'h00; 15'h5A2F: d <= 8'h7B;
                15'h5A30: d <= 8'h00; 15'h5A31: d <= 8'h00; 15'h5A32: d <= 8'h00; 15'h5A33: d <= 8'h00;
                15'h5A34: d <= 8'h00; 15'h5A35: d <= 8'h00; 15'h5A36: d <= 8'h00; 15'h5A37: d <= 8'h00;
                15'h5A38: d <= 8'h00; 15'h5A39: d <= 8'h00; 15'h5A3A: d <= 8'h00; 15'h5A3B: d <= 8'h00;
                15'h5A3C: d <= 8'h00; 15'h5A3D: d <= 8'h00; 15'h5A3E: d <= 8'h00; 15'h5A3F: d <= 8'h00;
                15'h5A40: d <= 8'h00; 15'h5A41: d <= 8'h00; 15'h5A42: d <= 8'h00; 15'h5A43: d <= 8'h00;
                15'h5A44: d <= 8'h00; 15'h5A45: d <= 8'h00; 15'h5A46: d <= 8'h00; 15'h5A47: d <= 8'h00;
                15'h5A48: d <= 8'h00; 15'h5A49: d <= 8'h00; 15'h5A4A: d <= 8'h00; 15'h5A4B: d <= 8'h00;
                15'h5A4C: d <= 8'h00; 15'h5A4D: d <= 8'h00; 15'h5A4E: d <= 8'h00; 15'h5A4F: d <= 8'h00;
                15'h5A50: d <= 8'h00; 15'h5A51: d <= 8'h00; 15'h5A52: d <= 8'h00; 15'h5A53: d <= 8'h00;
                15'h5A54: d <= 8'h00; 15'h5A55: d <= 8'h00; 15'h5A56: d <= 8'h00; 15'h5A57: d <= 8'h00;
                15'h5A58: d <= 8'h45; 15'h5A59: d <= 8'h35; 15'h5A5A: d <= 8'h32; 15'h5A5B: d <= 8'h00;
                15'h5A5C: d <= 8'h00; 15'h5A5D: d <= 8'h00; 15'h5A5E: d <= 8'h00; 15'h5A5F: d <= 8'h00;
                15'h5A60: d <= 8'h00; 15'h5A61: d <= 8'h00; 15'h5A62: d <= 8'h00; 15'h5A63: d <= 8'h00;
                15'h5A64: d <= 8'h00; 15'h5A65: d <= 8'h00; 15'h5A66: d <= 8'h00; 15'h5A67: d <= 8'h00;
                15'h5A68: d <= 8'h00; 15'h5A69: d <= 8'h00; 15'h5A6A: d <= 8'h00; 15'h5A6B: d <= 8'h00;
                15'h5A6C: d <= 8'h00; 15'h5A6D: d <= 8'h00; 15'h5A6E: d <= 8'h00; 15'h5A6F: d <= 8'h00;
                15'h5A70: d <= 8'h00; 15'h5A71: d <= 8'h00; 15'h5A72: d <= 8'h00; 15'h5A73: d <= 8'h00;
                15'h5A74: d <= 8'h00; 15'h5A75: d <= 8'h00; 15'h5A76: d <= 8'h00; 15'h5A77: d <= 8'h00;
                15'h5A78: d <= 8'h00; 15'h5A79: d <= 8'h00; 15'h5A7A: d <= 8'h00; 15'h5A7B: d <= 8'h00;
                15'h5A7C: d <= 8'h00; 15'h5A7D: d <= 8'h00; 15'h5A7E: d <= 8'h00; 15'h5A7F: d <= 8'hE0;
                15'h5A80: d <= 8'h10; 15'h5A81: d <= 8'h15; 15'h5A82: d <= 8'h1A; 15'h5A83: d <= 8'h1F;
                15'h5A84: d <= 8'h20; 15'h5A85: d <= 8'h25; 15'h5A86: d <= 8'h2A; 15'h5A87: d <= 8'h2F;
                15'h5A88: d <= 8'h34; 15'h5A89: d <= 8'h38; 15'h5A8A: d <= 8'h3C; 15'h5A8B: d <= 8'h31;
                15'h5A8C: d <= 8'h39; 15'h5A8D: d <= 8'h3D; 15'h5A8E: d <= 8'h32; 15'h5A8F: d <= 8'h36;
                15'h5A90: d <= 8'h3E; 15'h5A91: d <= 8'h33; 15'h5A92: d <= 8'h37; 15'h5A93: d <= 8'h3B;
                15'h5A94: d <= 8'h44; 15'h5A95: d <= 8'h48; 15'h5A96: d <= 8'h4C; 15'h5A97: d <= 8'h41;
                15'h5A98: d <= 8'h49; 15'h5A99: d <= 8'h4D; 15'h5A9A: d <= 8'h42; 15'h5A9B: d <= 8'h46;
                15'h5A9C: d <= 8'h4E; 15'h5A9D: d <= 8'h43; 15'h5A9E: d <= 8'h47; 15'h5A9F: d <= 8'h4B;
                15'h5AA0: d <= 8'h50; 15'h5AA1: d <= 8'h55; 15'h5AA2: d <= 8'h5A; 15'h5AA3: d <= 8'h5F;
                15'h5AA4: d <= 8'h60; 15'h5AA5: d <= 8'h65; 15'h5AA6: d <= 8'h6A; 15'h5AA7: d <= 8'h6F;
                15'h5AA8: d <= 8'h74; 15'h5AA9: d <= 8'h78; 15'h5AAA: d <= 8'h7C; 15'h5AAB: d <= 8'h71;
                15'h5AAC: d <= 8'h79; 15'h5AAD: d <= 8'h7D; 15'h5AAE: d <= 8'h72; 15'h5AAF: d <= 8'h76;
                15'h5AB0: d <= 8'h7E; 15'h5AB1: d <= 8'h73; 15'h5AB2: d <= 8'h77; 15'h5AB3: d <= 8'h7B;
                15'h5AB4: d <= 8'h84; 15'h5AB5: d <= 8'h88; 15'h5AB6: d <= 8'h8C; 15'h5AB7: d <= 8'h81;
                15'h5AB8: d <= 8'h89; 15'h5AB9: d <= 8'h8D; 15'h5ABA: d <= 8'h82; 15'h5ABB: d <= 8'h86;
                15'h5ABC: d <= 8'h8E; 15'h5ABD: d <= 8'h83; 15'h5ABE: d <= 8'h87; 15'h5ABF: d <= 8'h8B;
                15'h5AC0: d <= 8'h90; 15'h5AC1: d <= 8'h95; 15'h5AC2: d <= 8'h9A; 15'h5AC3: d <= 8'h9F;
                15'h5AC4: d <= 8'hA4; 15'h5AC5: d <= 8'hA8; 15'h5AC6: d <= 8'hAC; 15'h5AC7: d <= 8'hA1;
                15'h5AC8: d <= 8'hA9; 15'h5AC9: d <= 8'hAD; 15'h5ACA: d <= 8'hA2; 15'h5ACB: d <= 8'hA6;
                15'h5ACC: d <= 8'hAE; 15'h5ACD: d <= 8'hA3; 15'h5ACE: d <= 8'hA7; 15'h5ACF: d <= 8'hAB;
                15'h5AD0: d <= 8'hB4; 15'h5AD1: d <= 8'hB8; 15'h5AD2: d <= 8'hBC; 15'h5AD3: d <= 8'hB1;
                15'h5AD4: d <= 8'hB9; 15'h5AD5: d <= 8'hBD; 15'h5AD6: d <= 8'hB2; 15'h5AD7: d <= 8'hB6;
                15'h5AD8: d <= 8'hBE; 15'h5AD9: d <= 8'hB3; 15'h5ADA: d <= 8'hB7; 15'h5ADB: d <= 8'hBB;
                15'h5ADC: d <= 8'hC4; 15'h5ADD: d <= 8'hC8; 15'h5ADE: d <= 8'hCC; 15'h5ADF: d <= 8'hC1;
                15'h5AE0: d <= 8'hC9; 15'h5AE1: d <= 8'hCD; 15'h5AE2: d <= 8'hC2; 15'h5AE3: d <= 8'hC6;
                15'h5AE4: d <= 8'hCE; 15'h5AE5: d <= 8'hC3; 15'h5AE6: d <= 8'hC7; 15'h5AE7: d <= 8'hCB;
                15'h5AE8: d <= 8'hC0; 15'h5AE9: d <= 8'hC5; 15'h5AEA: d <= 8'hCA; 15'h5AEB: d <= 8'hCF;
                15'h5AEC: d <= 8'hD0; 15'h5AED: d <= 8'hD5; 15'h5AEE: d <= 8'hDA; 15'h5AEF: d <= 8'hDF;
                15'h5AF0: d <= 8'h74; 15'h5AF1: d <= 8'h78; 15'h5AF2: d <= 8'h7C; 15'h5AF3: d <= 8'h71;
                15'h5AF4: d <= 8'h79; 15'h5AF5: d <= 8'h7D; 15'h5AF6: d <= 8'h72; 15'h5AF7: d <= 8'h76;
                15'h5AF8: d <= 8'h7E; 15'h5AF9: d <= 8'h73; 15'h5AFA: d <= 8'h77; 15'h5AFB: d <= 8'h7B;
                15'h5AFC: d <= 8'hA0; 15'h5AFD: d <= 8'hA5; 15'h5AFE: d <= 8'hAA; 15'h5AFF: d <= 8'hAF;
                15'h5B00: d <= 8'h00; 15'h5B01: d <= 8'h00; 15'h5B02: d <= 8'h00; 15'h5B03: d <= 8'h00;
                15'h5B04: d <= 8'h00; 15'h5B05: d <= 8'h00; 15'h5B06: d <= 8'h00; 15'h5B07: d <= 8'h00;
                15'h5B08: d <= 8'h00; 15'h5B09: d <= 8'h00; 15'h5B0A: d <= 8'h00; 15'h5B0B: d <= 8'h00;
                15'h5B0C: d <= 8'h00; 15'h5B0D: d <= 8'h00; 15'h5B0E: d <= 8'h00; 15'h5B0F: d <= 8'h00;
                15'h5B10: d <= 8'h00; 15'h5B11: d <= 8'h00; 15'h5B12: d <= 8'h00; 15'h5B13: d <= 8'h00;
                15'h5B14: d <= 8'h00; 15'h5B15: d <= 8'h00; 15'h5B16: d <= 8'h00; 15'h5B17: d <= 8'h00;
                15'h5B18: d <= 8'h00; 15'h5B19: d <= 8'h00; 15'h5B1A: d <= 8'h00; 15'h5B1B: d <= 8'h00;
                15'h5B1C: d <= 8'h00; 15'h5B1D: d <= 8'h00; 15'h5B1E: d <= 8'h00; 15'h5B1F: d <= 8'h00;
                15'h5B20: d <= 8'h00; 15'h5B21: d <= 8'h00; 15'h5B22: d <= 8'h00; 15'h5B23: d <= 8'h00;
                15'h5B24: d <= 8'h00; 15'h5B25: d <= 8'h00; 15'h5B26: d <= 8'h00; 15'h5B27: d <= 8'h00;
                15'h5B28: d <= 8'h00; 15'h5B29: d <= 8'h00; 15'h5B2A: d <= 8'h00; 15'h5B2B: d <= 8'h00;
                15'h5B2C: d <= 8'h00; 15'h5B2D: d <= 8'h00; 15'h5B2E: d <= 8'h00; 15'h5B2F: d <= 8'h7B;
                15'h5B30: d <= 8'h00; 15'h5B31: d <= 8'h00; 15'h5B32: d <= 8'h00; 15'h5B33: d <= 8'h00;
                15'h5B34: d <= 8'h00; 15'h5B35: d <= 8'h00; 15'h5B36: d <= 8'h00; 15'h5B37: d <= 8'h00;
                15'h5B38: d <= 8'h00; 15'h5B39: d <= 8'h00; 15'h5B3A: d <= 8'h00; 15'h5B3B: d <= 8'h00;
                15'h5B3C: d <= 8'h00; 15'h5B3D: d <= 8'h00; 15'h5B3E: d <= 8'h00; 15'h5B3F: d <= 8'h00;
                15'h5B40: d <= 8'h00; 15'h5B41: d <= 8'h00; 15'h5B42: d <= 8'h00; 15'h5B43: d <= 8'h00;
                15'h5B44: d <= 8'h00; 15'h5B45: d <= 8'h00; 15'h5B46: d <= 8'h00; 15'h5B47: d <= 8'h00;
                15'h5B48: d <= 8'h00; 15'h5B49: d <= 8'h00; 15'h5B4A: d <= 8'h00; 15'h5B4B: d <= 8'h00;
                15'h5B4C: d <= 8'h00; 15'h5B4D: d <= 8'h00; 15'h5B4E: d <= 8'h00; 15'h5B4F: d <= 8'h00;
                15'h5B50: d <= 8'h00; 15'h5B51: d <= 8'h00; 15'h5B52: d <= 8'h00; 15'h5B53: d <= 8'h00;
                15'h5B54: d <= 8'h00; 15'h5B55: d <= 8'h00; 15'h5B56: d <= 8'h00; 15'h5B57: d <= 8'h00;
                15'h5B58: d <= 8'h45; 15'h5B59: d <= 8'h35; 15'h5B5A: d <= 8'h32; 15'h5B5B: d <= 8'h00;
                15'h5B5C: d <= 8'h00; 15'h5B5D: d <= 8'h00; 15'h5B5E: d <= 8'h00; 15'h5B5F: d <= 8'h00;
                15'h5B60: d <= 8'h00; 15'h5B61: d <= 8'h00; 15'h5B62: d <= 8'h00; 15'h5B63: d <= 8'h00;
                15'h5B64: d <= 8'h00; 15'h5B65: d <= 8'h00; 15'h5B66: d <= 8'h00; 15'h5B67: d <= 8'h00;
                15'h5B68: d <= 8'h00; 15'h5B69: d <= 8'h00; 15'h5B6A: d <= 8'h00; 15'h5B6B: d <= 8'h00;
                15'h5B6C: d <= 8'h00; 15'h5B6D: d <= 8'h00; 15'h5B6E: d <= 8'h00; 15'h5B6F: d <= 8'h00;
                15'h5B70: d <= 8'h00; 15'h5B71: d <= 8'h00; 15'h5B72: d <= 8'h00; 15'h5B73: d <= 8'h00;
                15'h5B74: d <= 8'h00; 15'h5B75: d <= 8'h00; 15'h5B76: d <= 8'h00; 15'h5B77: d <= 8'h00;
                15'h5B78: d <= 8'h00; 15'h5B79: d <= 8'h00; 15'h5B7A: d <= 8'h00; 15'h5B7B: d <= 8'h00;
                15'h5B7C: d <= 8'h00; 15'h5B7D: d <= 8'h00; 15'h5B7E: d <= 8'h00; 15'h5B7F: d <= 8'hE0;
                15'h5B80: d <= 8'h10; 15'h5B81: d <= 8'h15; 15'h5B82: d <= 8'h1A; 15'h5B83: d <= 8'h1F;
                15'h5B84: d <= 8'h20; 15'h5B85: d <= 8'h25; 15'h5B86: d <= 8'h2A; 15'h5B87: d <= 8'h2F;
                15'h5B88: d <= 8'h34; 15'h5B89: d <= 8'h38; 15'h5B8A: d <= 8'h3C; 15'h5B8B: d <= 8'h31;
                15'h5B8C: d <= 8'h39; 15'h5B8D: d <= 8'h3D; 15'h5B8E: d <= 8'h32; 15'h5B8F: d <= 8'h36;
                15'h5B90: d <= 8'h3E; 15'h5B91: d <= 8'h33; 15'h5B92: d <= 8'h37; 15'h5B93: d <= 8'h3B;
                15'h5B94: d <= 8'h44; 15'h5B95: d <= 8'h48; 15'h5B96: d <= 8'h4C; 15'h5B97: d <= 8'h41;
                15'h5B98: d <= 8'h49; 15'h5B99: d <= 8'h4D; 15'h5B9A: d <= 8'h42; 15'h5B9B: d <= 8'h46;
                15'h5B9C: d <= 8'h4E; 15'h5B9D: d <= 8'h43; 15'h5B9E: d <= 8'h47; 15'h5B9F: d <= 8'h4B;
                15'h5BA0: d <= 8'h50; 15'h5BA1: d <= 8'h55; 15'h5BA2: d <= 8'h5A; 15'h5BA3: d <= 8'h5F;
                15'h5BA4: d <= 8'h60; 15'h5BA5: d <= 8'h65; 15'h5BA6: d <= 8'h6A; 15'h5BA7: d <= 8'h6F;
                15'h5BA8: d <= 8'h74; 15'h5BA9: d <= 8'h78; 15'h5BAA: d <= 8'h7C; 15'h5BAB: d <= 8'h71;
                15'h5BAC: d <= 8'h79; 15'h5BAD: d <= 8'h7D; 15'h5BAE: d <= 8'h72; 15'h5BAF: d <= 8'h76;
                15'h5BB0: d <= 8'h7E; 15'h5BB1: d <= 8'h73; 15'h5BB2: d <= 8'h77; 15'h5BB3: d <= 8'h7B;
                15'h5BB4: d <= 8'h84; 15'h5BB5: d <= 8'h88; 15'h5BB6: d <= 8'h8C; 15'h5BB7: d <= 8'h81;
                15'h5BB8: d <= 8'h89; 15'h5BB9: d <= 8'h8D; 15'h5BBA: d <= 8'h82; 15'h5BBB: d <= 8'h86;
                15'h5BBC: d <= 8'h8E; 15'h5BBD: d <= 8'h83; 15'h5BBE: d <= 8'h87; 15'h5BBF: d <= 8'h8B;
                15'h5BC0: d <= 8'h90; 15'h5BC1: d <= 8'h95; 15'h5BC2: d <= 8'h9A; 15'h5BC3: d <= 8'h9F;
                15'h5BC4: d <= 8'hA4; 15'h5BC5: d <= 8'hA8; 15'h5BC6: d <= 8'hAC; 15'h5BC7: d <= 8'hA1;
                15'h5BC8: d <= 8'hA9; 15'h5BC9: d <= 8'hAD; 15'h5BCA: d <= 8'hA2; 15'h5BCB: d <= 8'hA6;
                15'h5BCC: d <= 8'hAE; 15'h5BCD: d <= 8'hA3; 15'h5BCE: d <= 8'hA7; 15'h5BCF: d <= 8'hAB;
                15'h5BD0: d <= 8'hB4; 15'h5BD1: d <= 8'hB8; 15'h5BD2: d <= 8'hBC; 15'h5BD3: d <= 8'hB1;
                15'h5BD4: d <= 8'hB9; 15'h5BD5: d <= 8'hBD; 15'h5BD6: d <= 8'hB2; 15'h5BD7: d <= 8'hB6;
                15'h5BD8: d <= 8'hBE; 15'h5BD9: d <= 8'hB3; 15'h5BDA: d <= 8'hB7; 15'h5BDB: d <= 8'hBB;
                15'h5BDC: d <= 8'hC4; 15'h5BDD: d <= 8'hC8; 15'h5BDE: d <= 8'hCC; 15'h5BDF: d <= 8'hC1;
                15'h5BE0: d <= 8'hC9; 15'h5BE1: d <= 8'hCD; 15'h5BE2: d <= 8'hC2; 15'h5BE3: d <= 8'hC6;
                15'h5BE4: d <= 8'hCE; 15'h5BE5: d <= 8'hC3; 15'h5BE6: d <= 8'hC7; 15'h5BE7: d <= 8'hCB;
                15'h5BE8: d <= 8'hC0; 15'h5BE9: d <= 8'hC5; 15'h5BEA: d <= 8'hCA; 15'h5BEB: d <= 8'hCF;
                15'h5BEC: d <= 8'hD0; 15'h5BED: d <= 8'hD5; 15'h5BEE: d <= 8'hDA; 15'h5BEF: d <= 8'hDF;
                15'h5BF0: d <= 8'h74; 15'h5BF1: d <= 8'h78; 15'h5BF2: d <= 8'h7C; 15'h5BF3: d <= 8'h71;
                15'h5BF4: d <= 8'h79; 15'h5BF5: d <= 8'h7D; 15'h5BF6: d <= 8'h72; 15'h5BF7: d <= 8'h76;
                15'h5BF8: d <= 8'h7E; 15'h5BF9: d <= 8'h73; 15'h5BFA: d <= 8'h77; 15'h5BFB: d <= 8'h7B;
                15'h5BFC: d <= 8'hA0; 15'h5BFD: d <= 8'hA5; 15'h5BFE: d <= 8'hAA; 15'h5BFF: d <= 8'hAF;
                15'h5C00: d <= 8'h00; 15'h5C01: d <= 8'h00; 15'h5C02: d <= 8'h00; 15'h5C03: d <= 8'h00;
                15'h5C04: d <= 8'h00; 15'h5C05: d <= 8'h00; 15'h5C06: d <= 8'h00; 15'h5C07: d <= 8'h00;
                15'h5C08: d <= 8'h00; 15'h5C09: d <= 8'h00; 15'h5C0A: d <= 8'h00; 15'h5C0B: d <= 8'h00;
                15'h5C0C: d <= 8'h00; 15'h5C0D: d <= 8'h00; 15'h5C0E: d <= 8'h00; 15'h5C0F: d <= 8'h00;
                15'h5C10: d <= 8'h00; 15'h5C11: d <= 8'h00; 15'h5C12: d <= 8'h00; 15'h5C13: d <= 8'h00;
                15'h5C14: d <= 8'h00; 15'h5C15: d <= 8'h00; 15'h5C16: d <= 8'h00; 15'h5C17: d <= 8'h00;
                15'h5C18: d <= 8'h00; 15'h5C19: d <= 8'h00; 15'h5C1A: d <= 8'h00; 15'h5C1B: d <= 8'h00;
                15'h5C1C: d <= 8'h00; 15'h5C1D: d <= 8'h00; 15'h5C1E: d <= 8'h00; 15'h5C1F: d <= 8'h00;
                15'h5C20: d <= 8'h00; 15'h5C21: d <= 8'h00; 15'h5C22: d <= 8'h00; 15'h5C23: d <= 8'h00;
                15'h5C24: d <= 8'h00; 15'h5C25: d <= 8'h00; 15'h5C26: d <= 8'h00; 15'h5C27: d <= 8'h00;
                15'h5C28: d <= 8'h00; 15'h5C29: d <= 8'h00; 15'h5C2A: d <= 8'h00; 15'h5C2B: d <= 8'h00;
                15'h5C2C: d <= 8'h00; 15'h5C2D: d <= 8'h00; 15'h5C2E: d <= 8'h00; 15'h5C2F: d <= 8'h7B;
                15'h5C30: d <= 8'h00; 15'h5C31: d <= 8'h00; 15'h5C32: d <= 8'h00; 15'h5C33: d <= 8'h00;
                15'h5C34: d <= 8'h00; 15'h5C35: d <= 8'h00; 15'h5C36: d <= 8'h00; 15'h5C37: d <= 8'h00;
                15'h5C38: d <= 8'h00; 15'h5C39: d <= 8'h00; 15'h5C3A: d <= 8'h00; 15'h5C3B: d <= 8'h00;
                15'h5C3C: d <= 8'h00; 15'h5C3D: d <= 8'h00; 15'h5C3E: d <= 8'h00; 15'h5C3F: d <= 8'h00;
                15'h5C40: d <= 8'h00; 15'h5C41: d <= 8'h00; 15'h5C42: d <= 8'h00; 15'h5C43: d <= 8'h00;
                15'h5C44: d <= 8'h00; 15'h5C45: d <= 8'h00; 15'h5C46: d <= 8'h00; 15'h5C47: d <= 8'h00;
                15'h5C48: d <= 8'h00; 15'h5C49: d <= 8'h00; 15'h5C4A: d <= 8'h00; 15'h5C4B: d <= 8'h00;
                15'h5C4C: d <= 8'h00; 15'h5C4D: d <= 8'h00; 15'h5C4E: d <= 8'h00; 15'h5C4F: d <= 8'h00;
                15'h5C50: d <= 8'h00; 15'h5C51: d <= 8'h00; 15'h5C52: d <= 8'h00; 15'h5C53: d <= 8'h00;
                15'h5C54: d <= 8'h00; 15'h5C55: d <= 8'h00; 15'h5C56: d <= 8'h00; 15'h5C57: d <= 8'h00;
                15'h5C58: d <= 8'h45; 15'h5C59: d <= 8'h35; 15'h5C5A: d <= 8'h32; 15'h5C5B: d <= 8'h00;
                15'h5C5C: d <= 8'h00; 15'h5C5D: d <= 8'h00; 15'h5C5E: d <= 8'h00; 15'h5C5F: d <= 8'h00;
                15'h5C60: d <= 8'h00; 15'h5C61: d <= 8'h00; 15'h5C62: d <= 8'h00; 15'h5C63: d <= 8'h00;
                15'h5C64: d <= 8'h00; 15'h5C65: d <= 8'h00; 15'h5C66: d <= 8'h00; 15'h5C67: d <= 8'h00;
                15'h5C68: d <= 8'h00; 15'h5C69: d <= 8'h00; 15'h5C6A: d <= 8'h00; 15'h5C6B: d <= 8'h00;
                15'h5C6C: d <= 8'h00; 15'h5C6D: d <= 8'h00; 15'h5C6E: d <= 8'h00; 15'h5C6F: d <= 8'h00;
                15'h5C70: d <= 8'h00; 15'h5C71: d <= 8'h00; 15'h5C72: d <= 8'h00; 15'h5C73: d <= 8'h00;
                15'h5C74: d <= 8'h00; 15'h5C75: d <= 8'h00; 15'h5C76: d <= 8'h00; 15'h5C77: d <= 8'h00;
                15'h5C78: d <= 8'h00; 15'h5C79: d <= 8'h00; 15'h5C7A: d <= 8'h00; 15'h5C7B: d <= 8'h00;
                15'h5C7C: d <= 8'h00; 15'h5C7D: d <= 8'h00; 15'h5C7E: d <= 8'h00; 15'h5C7F: d <= 8'hE0;
                15'h5C80: d <= 8'h10; 15'h5C81: d <= 8'h15; 15'h5C82: d <= 8'h1A; 15'h5C83: d <= 8'h1F;
                15'h5C84: d <= 8'h20; 15'h5C85: d <= 8'h25; 15'h5C86: d <= 8'h2A; 15'h5C87: d <= 8'h2F;
                15'h5C88: d <= 8'h34; 15'h5C89: d <= 8'h38; 15'h5C8A: d <= 8'h3C; 15'h5C8B: d <= 8'h31;
                15'h5C8C: d <= 8'h39; 15'h5C8D: d <= 8'h3D; 15'h5C8E: d <= 8'h32; 15'h5C8F: d <= 8'h36;
                15'h5C90: d <= 8'h3E; 15'h5C91: d <= 8'h33; 15'h5C92: d <= 8'h37; 15'h5C93: d <= 8'h3B;
                15'h5C94: d <= 8'h44; 15'h5C95: d <= 8'h48; 15'h5C96: d <= 8'h4C; 15'h5C97: d <= 8'h41;
                15'h5C98: d <= 8'h49; 15'h5C99: d <= 8'h4D; 15'h5C9A: d <= 8'h42; 15'h5C9B: d <= 8'h46;
                15'h5C9C: d <= 8'h4E; 15'h5C9D: d <= 8'h43; 15'h5C9E: d <= 8'h47; 15'h5C9F: d <= 8'h4B;
                15'h5CA0: d <= 8'h50; 15'h5CA1: d <= 8'h55; 15'h5CA2: d <= 8'h5A; 15'h5CA3: d <= 8'h5F;
                15'h5CA4: d <= 8'h60; 15'h5CA5: d <= 8'h65; 15'h5CA6: d <= 8'h6A; 15'h5CA7: d <= 8'h6F;
                15'h5CA8: d <= 8'h74; 15'h5CA9: d <= 8'h78; 15'h5CAA: d <= 8'h7C; 15'h5CAB: d <= 8'h71;
                15'h5CAC: d <= 8'h79; 15'h5CAD: d <= 8'h7D; 15'h5CAE: d <= 8'h72; 15'h5CAF: d <= 8'h76;
                15'h5CB0: d <= 8'h7E; 15'h5CB1: d <= 8'h73; 15'h5CB2: d <= 8'h77; 15'h5CB3: d <= 8'h7B;
                15'h5CB4: d <= 8'h84; 15'h5CB5: d <= 8'h88; 15'h5CB6: d <= 8'h8C; 15'h5CB7: d <= 8'h81;
                15'h5CB8: d <= 8'h89; 15'h5CB9: d <= 8'h8D; 15'h5CBA: d <= 8'h82; 15'h5CBB: d <= 8'h86;
                15'h5CBC: d <= 8'h8E; 15'h5CBD: d <= 8'h83; 15'h5CBE: d <= 8'h87; 15'h5CBF: d <= 8'h8B;
                15'h5CC0: d <= 8'h90; 15'h5CC1: d <= 8'h95; 15'h5CC2: d <= 8'h9A; 15'h5CC3: d <= 8'h9F;
                15'h5CC4: d <= 8'hA4; 15'h5CC5: d <= 8'hA8; 15'h5CC6: d <= 8'hAC; 15'h5CC7: d <= 8'hA1;
                15'h5CC8: d <= 8'hA9; 15'h5CC9: d <= 8'hAD; 15'h5CCA: d <= 8'hA2; 15'h5CCB: d <= 8'hA6;
                15'h5CCC: d <= 8'hAE; 15'h5CCD: d <= 8'hA3; 15'h5CCE: d <= 8'hA7; 15'h5CCF: d <= 8'hAB;
                15'h5CD0: d <= 8'hB4; 15'h5CD1: d <= 8'hB8; 15'h5CD2: d <= 8'hBC; 15'h5CD3: d <= 8'hB1;
                15'h5CD4: d <= 8'hB9; 15'h5CD5: d <= 8'hBD; 15'h5CD6: d <= 8'hB2; 15'h5CD7: d <= 8'hB6;
                15'h5CD8: d <= 8'hBE; 15'h5CD9: d <= 8'hB3; 15'h5CDA: d <= 8'hB7; 15'h5CDB: d <= 8'hBB;
                15'h5CDC: d <= 8'hC4; 15'h5CDD: d <= 8'hC8; 15'h5CDE: d <= 8'hCC; 15'h5CDF: d <= 8'hC1;
                15'h5CE0: d <= 8'hC9; 15'h5CE1: d <= 8'hCD; 15'h5CE2: d <= 8'hC2; 15'h5CE3: d <= 8'hC6;
                15'h5CE4: d <= 8'hCE; 15'h5CE5: d <= 8'hC3; 15'h5CE6: d <= 8'hC7; 15'h5CE7: d <= 8'hCB;
                15'h5CE8: d <= 8'hC0; 15'h5CE9: d <= 8'hC5; 15'h5CEA: d <= 8'hCA; 15'h5CEB: d <= 8'hCF;
                15'h5CEC: d <= 8'hD0; 15'h5CED: d <= 8'hD5; 15'h5CEE: d <= 8'hDA; 15'h5CEF: d <= 8'hDF;
                15'h5CF0: d <= 8'h74; 15'h5CF1: d <= 8'h78; 15'h5CF2: d <= 8'h7C; 15'h5CF3: d <= 8'h71;
                15'h5CF4: d <= 8'h79; 15'h5CF5: d <= 8'h7D; 15'h5CF6: d <= 8'h72; 15'h5CF7: d <= 8'h76;
                15'h5CF8: d <= 8'h7E; 15'h5CF9: d <= 8'h73; 15'h5CFA: d <= 8'h77; 15'h5CFB: d <= 8'h7B;
                15'h5CFC: d <= 8'hA0; 15'h5CFD: d <= 8'hA5; 15'h5CFE: d <= 8'hAA; 15'h5CFF: d <= 8'hAF;
                15'h5D00: d <= 8'h00; 15'h5D01: d <= 8'h00; 15'h5D02: d <= 8'h00; 15'h5D03: d <= 8'h00;
                15'h5D04: d <= 8'h00; 15'h5D05: d <= 8'h00; 15'h5D06: d <= 8'h00; 15'h5D07: d <= 8'h00;
                15'h5D08: d <= 8'h00; 15'h5D09: d <= 8'h00; 15'h5D0A: d <= 8'h00; 15'h5D0B: d <= 8'h00;
                15'h5D0C: d <= 8'h00; 15'h5D0D: d <= 8'h00; 15'h5D0E: d <= 8'h00; 15'h5D0F: d <= 8'h00;
                15'h5D10: d <= 8'h00; 15'h5D11: d <= 8'h00; 15'h5D12: d <= 8'h00; 15'h5D13: d <= 8'h00;
                15'h5D14: d <= 8'h00; 15'h5D15: d <= 8'h00; 15'h5D16: d <= 8'h00; 15'h5D17: d <= 8'h00;
                15'h5D18: d <= 8'h00; 15'h5D19: d <= 8'h00; 15'h5D1A: d <= 8'h00; 15'h5D1B: d <= 8'h00;
                15'h5D1C: d <= 8'h00; 15'h5D1D: d <= 8'h00; 15'h5D1E: d <= 8'h00; 15'h5D1F: d <= 8'h00;
                15'h5D20: d <= 8'h00; 15'h5D21: d <= 8'h00; 15'h5D22: d <= 8'h00; 15'h5D23: d <= 8'h00;
                15'h5D24: d <= 8'h00; 15'h5D25: d <= 8'h00; 15'h5D26: d <= 8'h00; 15'h5D27: d <= 8'h00;
                15'h5D28: d <= 8'h00; 15'h5D29: d <= 8'h00; 15'h5D2A: d <= 8'h00; 15'h5D2B: d <= 8'h00;
                15'h5D2C: d <= 8'h00; 15'h5D2D: d <= 8'h00; 15'h5D2E: d <= 8'h00; 15'h5D2F: d <= 8'h7B;
                15'h5D30: d <= 8'h00; 15'h5D31: d <= 8'h00; 15'h5D32: d <= 8'h00; 15'h5D33: d <= 8'h00;
                15'h5D34: d <= 8'h00; 15'h5D35: d <= 8'h00; 15'h5D36: d <= 8'h00; 15'h5D37: d <= 8'h00;
                15'h5D38: d <= 8'h00; 15'h5D39: d <= 8'h00; 15'h5D3A: d <= 8'h00; 15'h5D3B: d <= 8'h00;
                15'h5D3C: d <= 8'h00; 15'h5D3D: d <= 8'h00; 15'h5D3E: d <= 8'h00; 15'h5D3F: d <= 8'h00;
                15'h5D40: d <= 8'h00; 15'h5D41: d <= 8'h00; 15'h5D42: d <= 8'h00; 15'h5D43: d <= 8'h00;
                15'h5D44: d <= 8'h00; 15'h5D45: d <= 8'h00; 15'h5D46: d <= 8'h00; 15'h5D47: d <= 8'h00;
                15'h5D48: d <= 8'h00; 15'h5D49: d <= 8'h00; 15'h5D4A: d <= 8'h00; 15'h5D4B: d <= 8'h00;
                15'h5D4C: d <= 8'h00; 15'h5D4D: d <= 8'h00; 15'h5D4E: d <= 8'h00; 15'h5D4F: d <= 8'h00;
                15'h5D50: d <= 8'h00; 15'h5D51: d <= 8'h00; 15'h5D52: d <= 8'h00; 15'h5D53: d <= 8'h00;
                15'h5D54: d <= 8'h00; 15'h5D55: d <= 8'h00; 15'h5D56: d <= 8'h00; 15'h5D57: d <= 8'h00;
                15'h5D58: d <= 8'h45; 15'h5D59: d <= 8'h35; 15'h5D5A: d <= 8'h32; 15'h5D5B: d <= 8'h00;
                15'h5D5C: d <= 8'h00; 15'h5D5D: d <= 8'h00; 15'h5D5E: d <= 8'h00; 15'h5D5F: d <= 8'h00;
                15'h5D60: d <= 8'h00; 15'h5D61: d <= 8'h00; 15'h5D62: d <= 8'h00; 15'h5D63: d <= 8'h00;
                15'h5D64: d <= 8'h00; 15'h5D65: d <= 8'h00; 15'h5D66: d <= 8'h00; 15'h5D67: d <= 8'h00;
                15'h5D68: d <= 8'h00; 15'h5D69: d <= 8'h00; 15'h5D6A: d <= 8'h00; 15'h5D6B: d <= 8'h00;
                15'h5D6C: d <= 8'h00; 15'h5D6D: d <= 8'h00; 15'h5D6E: d <= 8'h00; 15'h5D6F: d <= 8'h00;
                15'h5D70: d <= 8'h00; 15'h5D71: d <= 8'h00; 15'h5D72: d <= 8'h00; 15'h5D73: d <= 8'h00;
                15'h5D74: d <= 8'h00; 15'h5D75: d <= 8'h00; 15'h5D76: d <= 8'h00; 15'h5D77: d <= 8'h00;
                15'h5D78: d <= 8'h00; 15'h5D79: d <= 8'h00; 15'h5D7A: d <= 8'h00; 15'h5D7B: d <= 8'h00;
                15'h5D7C: d <= 8'h00; 15'h5D7D: d <= 8'h00; 15'h5D7E: d <= 8'h00; 15'h5D7F: d <= 8'hE0;
                15'h5D80: d <= 8'h10; 15'h5D81: d <= 8'h15; 15'h5D82: d <= 8'h1A; 15'h5D83: d <= 8'h1F;
                15'h5D84: d <= 8'h20; 15'h5D85: d <= 8'h25; 15'h5D86: d <= 8'h2A; 15'h5D87: d <= 8'h2F;
                15'h5D88: d <= 8'h34; 15'h5D89: d <= 8'h38; 15'h5D8A: d <= 8'h3C; 15'h5D8B: d <= 8'h31;
                15'h5D8C: d <= 8'h39; 15'h5D8D: d <= 8'h3D; 15'h5D8E: d <= 8'h32; 15'h5D8F: d <= 8'h36;
                15'h5D90: d <= 8'h3E; 15'h5D91: d <= 8'h33; 15'h5D92: d <= 8'h37; 15'h5D93: d <= 8'h3B;
                15'h5D94: d <= 8'h44; 15'h5D95: d <= 8'h48; 15'h5D96: d <= 8'h4C; 15'h5D97: d <= 8'h41;
                15'h5D98: d <= 8'h49; 15'h5D99: d <= 8'h4D; 15'h5D9A: d <= 8'h42; 15'h5D9B: d <= 8'h46;
                15'h5D9C: d <= 8'h4E; 15'h5D9D: d <= 8'h43; 15'h5D9E: d <= 8'h47; 15'h5D9F: d <= 8'h4B;
                15'h5DA0: d <= 8'h50; 15'h5DA1: d <= 8'h55; 15'h5DA2: d <= 8'h5A; 15'h5DA3: d <= 8'h5F;
                15'h5DA4: d <= 8'h60; 15'h5DA5: d <= 8'h65; 15'h5DA6: d <= 8'h6A; 15'h5DA7: d <= 8'h6F;
                15'h5DA8: d <= 8'h74; 15'h5DA9: d <= 8'h78; 15'h5DAA: d <= 8'h7C; 15'h5DAB: d <= 8'h71;
                15'h5DAC: d <= 8'h79; 15'h5DAD: d <= 8'h7D; 15'h5DAE: d <= 8'h72; 15'h5DAF: d <= 8'h76;
                15'h5DB0: d <= 8'h7E; 15'h5DB1: d <= 8'h73; 15'h5DB2: d <= 8'h77; 15'h5DB3: d <= 8'h7B;
                15'h5DB4: d <= 8'h84; 15'h5DB5: d <= 8'h88; 15'h5DB6: d <= 8'h8C; 15'h5DB7: d <= 8'h81;
                15'h5DB8: d <= 8'h89; 15'h5DB9: d <= 8'h8D; 15'h5DBA: d <= 8'h82; 15'h5DBB: d <= 8'h86;
                15'h5DBC: d <= 8'h8E; 15'h5DBD: d <= 8'h83; 15'h5DBE: d <= 8'h87; 15'h5DBF: d <= 8'h8B;
                15'h5DC0: d <= 8'h90; 15'h5DC1: d <= 8'h95; 15'h5DC2: d <= 8'h9A; 15'h5DC3: d <= 8'h9F;
                15'h5DC4: d <= 8'hA4; 15'h5DC5: d <= 8'hA8; 15'h5DC6: d <= 8'hAC; 15'h5DC7: d <= 8'hA1;
                15'h5DC8: d <= 8'hA9; 15'h5DC9: d <= 8'hAD; 15'h5DCA: d <= 8'hA2; 15'h5DCB: d <= 8'hA6;
                15'h5DCC: d <= 8'hAE; 15'h5DCD: d <= 8'hA3; 15'h5DCE: d <= 8'hA7; 15'h5DCF: d <= 8'hAB;
                15'h5DD0: d <= 8'hB4; 15'h5DD1: d <= 8'hB8; 15'h5DD2: d <= 8'hBC; 15'h5DD3: d <= 8'hB1;
                15'h5DD4: d <= 8'hB9; 15'h5DD5: d <= 8'hBD; 15'h5DD6: d <= 8'hB2; 15'h5DD7: d <= 8'hB6;
                15'h5DD8: d <= 8'hBE; 15'h5DD9: d <= 8'hB3; 15'h5DDA: d <= 8'hB7; 15'h5DDB: d <= 8'hBB;
                15'h5DDC: d <= 8'hC4; 15'h5DDD: d <= 8'hC8; 15'h5DDE: d <= 8'hCC; 15'h5DDF: d <= 8'hC1;
                15'h5DE0: d <= 8'hC9; 15'h5DE1: d <= 8'hCD; 15'h5DE2: d <= 8'hC2; 15'h5DE3: d <= 8'hC6;
                15'h5DE4: d <= 8'hCE; 15'h5DE5: d <= 8'hC3; 15'h5DE6: d <= 8'hC7; 15'h5DE7: d <= 8'hCB;
                15'h5DE8: d <= 8'hC0; 15'h5DE9: d <= 8'hC5; 15'h5DEA: d <= 8'hCA; 15'h5DEB: d <= 8'hCF;
                15'h5DEC: d <= 8'hD0; 15'h5DED: d <= 8'hD5; 15'h5DEE: d <= 8'hDA; 15'h5DEF: d <= 8'hDF;
                15'h5DF0: d <= 8'h74; 15'h5DF1: d <= 8'h78; 15'h5DF2: d <= 8'h7C; 15'h5DF3: d <= 8'h71;
                15'h5DF4: d <= 8'h79; 15'h5DF5: d <= 8'h7D; 15'h5DF6: d <= 8'h72; 15'h5DF7: d <= 8'h76;
                15'h5DF8: d <= 8'h7E; 15'h5DF9: d <= 8'h73; 15'h5DFA: d <= 8'h77; 15'h5DFB: d <= 8'h7B;
                15'h5DFC: d <= 8'hA0; 15'h5DFD: d <= 8'hA5; 15'h5DFE: d <= 8'hAA; 15'h5DFF: d <= 8'hAF;
                15'h5E00: d <= 8'h00; 15'h5E01: d <= 8'h00; 15'h5E02: d <= 8'h00; 15'h5E03: d <= 8'h00;
                15'h5E04: d <= 8'h00; 15'h5E05: d <= 8'h00; 15'h5E06: d <= 8'h00; 15'h5E07: d <= 8'h00;
                15'h5E08: d <= 8'h00; 15'h5E09: d <= 8'h00; 15'h5E0A: d <= 8'h00; 15'h5E0B: d <= 8'h00;
                15'h5E0C: d <= 8'h00; 15'h5E0D: d <= 8'h00; 15'h5E0E: d <= 8'h00; 15'h5E0F: d <= 8'h00;
                15'h5E10: d <= 8'h00; 15'h5E11: d <= 8'h00; 15'h5E12: d <= 8'h00; 15'h5E13: d <= 8'h00;
                15'h5E14: d <= 8'h00; 15'h5E15: d <= 8'h00; 15'h5E16: d <= 8'h00; 15'h5E17: d <= 8'h00;
                15'h5E18: d <= 8'h00; 15'h5E19: d <= 8'h00; 15'h5E1A: d <= 8'h00; 15'h5E1B: d <= 8'h00;
                15'h5E1C: d <= 8'h00; 15'h5E1D: d <= 8'h00; 15'h5E1E: d <= 8'h00; 15'h5E1F: d <= 8'h00;
                15'h5E20: d <= 8'h00; 15'h5E21: d <= 8'h00; 15'h5E22: d <= 8'h00; 15'h5E23: d <= 8'h00;
                15'h5E24: d <= 8'h00; 15'h5E25: d <= 8'h00; 15'h5E26: d <= 8'h00; 15'h5E27: d <= 8'h00;
                15'h5E28: d <= 8'h00; 15'h5E29: d <= 8'h00; 15'h5E2A: d <= 8'h00; 15'h5E2B: d <= 8'h00;
                15'h5E2C: d <= 8'h00; 15'h5E2D: d <= 8'h00; 15'h5E2E: d <= 8'h00; 15'h5E2F: d <= 8'h7B;
                15'h5E30: d <= 8'h00; 15'h5E31: d <= 8'h00; 15'h5E32: d <= 8'h00; 15'h5E33: d <= 8'h00;
                15'h5E34: d <= 8'h00; 15'h5E35: d <= 8'h00; 15'h5E36: d <= 8'h00; 15'h5E37: d <= 8'h00;
                15'h5E38: d <= 8'h00; 15'h5E39: d <= 8'h00; 15'h5E3A: d <= 8'h00; 15'h5E3B: d <= 8'h00;
                15'h5E3C: d <= 8'h00; 15'h5E3D: d <= 8'h00; 15'h5E3E: d <= 8'h00; 15'h5E3F: d <= 8'h00;
                15'h5E40: d <= 8'h00; 15'h5E41: d <= 8'h00; 15'h5E42: d <= 8'h00; 15'h5E43: d <= 8'h00;
                15'h5E44: d <= 8'h00; 15'h5E45: d <= 8'h00; 15'h5E46: d <= 8'h00; 15'h5E47: d <= 8'h00;
                15'h5E48: d <= 8'h00; 15'h5E49: d <= 8'h00; 15'h5E4A: d <= 8'h00; 15'h5E4B: d <= 8'h00;
                15'h5E4C: d <= 8'h00; 15'h5E4D: d <= 8'h00; 15'h5E4E: d <= 8'h00; 15'h5E4F: d <= 8'h00;
                15'h5E50: d <= 8'h00; 15'h5E51: d <= 8'h00; 15'h5E52: d <= 8'h00; 15'h5E53: d <= 8'h00;
                15'h5E54: d <= 8'h00; 15'h5E55: d <= 8'h00; 15'h5E56: d <= 8'h00; 15'h5E57: d <= 8'h00;
                15'h5E58: d <= 8'h45; 15'h5E59: d <= 8'h35; 15'h5E5A: d <= 8'h32; 15'h5E5B: d <= 8'h00;
                15'h5E5C: d <= 8'h00; 15'h5E5D: d <= 8'h00; 15'h5E5E: d <= 8'h00; 15'h5E5F: d <= 8'h00;
                15'h5E60: d <= 8'h00; 15'h5E61: d <= 8'h00; 15'h5E62: d <= 8'h00; 15'h5E63: d <= 8'h00;
                15'h5E64: d <= 8'h00; 15'h5E65: d <= 8'h00; 15'h5E66: d <= 8'h00; 15'h5E67: d <= 8'h00;
                15'h5E68: d <= 8'h00; 15'h5E69: d <= 8'h00; 15'h5E6A: d <= 8'h00; 15'h5E6B: d <= 8'h00;
                15'h5E6C: d <= 8'h00; 15'h5E6D: d <= 8'h00; 15'h5E6E: d <= 8'h00; 15'h5E6F: d <= 8'h00;
                15'h5E70: d <= 8'h00; 15'h5E71: d <= 8'h00; 15'h5E72: d <= 8'h00; 15'h5E73: d <= 8'h00;
                15'h5E74: d <= 8'h00; 15'h5E75: d <= 8'h00; 15'h5E76: d <= 8'h00; 15'h5E77: d <= 8'h00;
                15'h5E78: d <= 8'h00; 15'h5E79: d <= 8'h00; 15'h5E7A: d <= 8'h00; 15'h5E7B: d <= 8'h00;
                15'h5E7C: d <= 8'h00; 15'h5E7D: d <= 8'h00; 15'h5E7E: d <= 8'h00; 15'h5E7F: d <= 8'hE0;
                15'h5E80: d <= 8'h10; 15'h5E81: d <= 8'h15; 15'h5E82: d <= 8'h1A; 15'h5E83: d <= 8'h1F;
                15'h5E84: d <= 8'h20; 15'h5E85: d <= 8'h25; 15'h5E86: d <= 8'h2A; 15'h5E87: d <= 8'h2F;
                15'h5E88: d <= 8'h34; 15'h5E89: d <= 8'h38; 15'h5E8A: d <= 8'h3C; 15'h5E8B: d <= 8'h31;
                15'h5E8C: d <= 8'h39; 15'h5E8D: d <= 8'h3D; 15'h5E8E: d <= 8'h32; 15'h5E8F: d <= 8'h36;
                15'h5E90: d <= 8'h3E; 15'h5E91: d <= 8'h33; 15'h5E92: d <= 8'h37; 15'h5E93: d <= 8'h3B;
                15'h5E94: d <= 8'h44; 15'h5E95: d <= 8'h48; 15'h5E96: d <= 8'h4C; 15'h5E97: d <= 8'h41;
                15'h5E98: d <= 8'h49; 15'h5E99: d <= 8'h4D; 15'h5E9A: d <= 8'h42; 15'h5E9B: d <= 8'h46;
                15'h5E9C: d <= 8'h4E; 15'h5E9D: d <= 8'h43; 15'h5E9E: d <= 8'h47; 15'h5E9F: d <= 8'h4B;
                15'h5EA0: d <= 8'h50; 15'h5EA1: d <= 8'h55; 15'h5EA2: d <= 8'h5A; 15'h5EA3: d <= 8'h5F;
                15'h5EA4: d <= 8'h60; 15'h5EA5: d <= 8'h65; 15'h5EA6: d <= 8'h6A; 15'h5EA7: d <= 8'h6F;
                15'h5EA8: d <= 8'h74; 15'h5EA9: d <= 8'h78; 15'h5EAA: d <= 8'h7C; 15'h5EAB: d <= 8'h71;
                15'h5EAC: d <= 8'h79; 15'h5EAD: d <= 8'h7D; 15'h5EAE: d <= 8'h72; 15'h5EAF: d <= 8'h76;
                15'h5EB0: d <= 8'h7E; 15'h5EB1: d <= 8'h73; 15'h5EB2: d <= 8'h77; 15'h5EB3: d <= 8'h7B;
                15'h5EB4: d <= 8'h84; 15'h5EB5: d <= 8'h88; 15'h5EB6: d <= 8'h8C; 15'h5EB7: d <= 8'h81;
                15'h5EB8: d <= 8'h89; 15'h5EB9: d <= 8'h8D; 15'h5EBA: d <= 8'h82; 15'h5EBB: d <= 8'h86;
                15'h5EBC: d <= 8'h8E; 15'h5EBD: d <= 8'h83; 15'h5EBE: d <= 8'h87; 15'h5EBF: d <= 8'h8B;
                15'h5EC0: d <= 8'h90; 15'h5EC1: d <= 8'h95; 15'h5EC2: d <= 8'h9A; 15'h5EC3: d <= 8'h9F;
                15'h5EC4: d <= 8'hA4; 15'h5EC5: d <= 8'hA8; 15'h5EC6: d <= 8'hAC; 15'h5EC7: d <= 8'hA1;
                15'h5EC8: d <= 8'hA9; 15'h5EC9: d <= 8'hAD; 15'h5ECA: d <= 8'hA2; 15'h5ECB: d <= 8'hA6;
                15'h5ECC: d <= 8'hAE; 15'h5ECD: d <= 8'hA3; 15'h5ECE: d <= 8'hA7; 15'h5ECF: d <= 8'hAB;
                15'h5ED0: d <= 8'hB4; 15'h5ED1: d <= 8'hB8; 15'h5ED2: d <= 8'hBC; 15'h5ED3: d <= 8'hB1;
                15'h5ED4: d <= 8'hB9; 15'h5ED5: d <= 8'hBD; 15'h5ED6: d <= 8'hB2; 15'h5ED7: d <= 8'hB6;
                15'h5ED8: d <= 8'hBE; 15'h5ED9: d <= 8'hB3; 15'h5EDA: d <= 8'hB7; 15'h5EDB: d <= 8'hBB;
                15'h5EDC: d <= 8'hC4; 15'h5EDD: d <= 8'hC8; 15'h5EDE: d <= 8'hCC; 15'h5EDF: d <= 8'hC1;
                15'h5EE0: d <= 8'hC9; 15'h5EE1: d <= 8'hCD; 15'h5EE2: d <= 8'hC2; 15'h5EE3: d <= 8'hC6;
                15'h5EE4: d <= 8'hCE; 15'h5EE5: d <= 8'hC3; 15'h5EE6: d <= 8'hC7; 15'h5EE7: d <= 8'hCB;
                15'h5EE8: d <= 8'hC0; 15'h5EE9: d <= 8'hC5; 15'h5EEA: d <= 8'hCA; 15'h5EEB: d <= 8'hCF;
                15'h5EEC: d <= 8'hD0; 15'h5EED: d <= 8'hD5; 15'h5EEE: d <= 8'hDA; 15'h5EEF: d <= 8'hDF;
                15'h5EF0: d <= 8'h74; 15'h5EF1: d <= 8'h78; 15'h5EF2: d <= 8'h7C; 15'h5EF3: d <= 8'h71;
                15'h5EF4: d <= 8'h79; 15'h5EF5: d <= 8'h7D; 15'h5EF6: d <= 8'h72; 15'h5EF7: d <= 8'h76;
                15'h5EF8: d <= 8'h7E; 15'h5EF9: d <= 8'h73; 15'h5EFA: d <= 8'h77; 15'h5EFB: d <= 8'h7B;
                15'h5EFC: d <= 8'hA0; 15'h5EFD: d <= 8'hA5; 15'h5EFE: d <= 8'hAA; 15'h5EFF: d <= 8'hAF;
                15'h5F00: d <= 8'h00; 15'h5F01: d <= 8'h00; 15'h5F02: d <= 8'h00; 15'h5F03: d <= 8'h00;
                15'h5F04: d <= 8'h00; 15'h5F05: d <= 8'h00; 15'h5F06: d <= 8'h00; 15'h5F07: d <= 8'h00;
                15'h5F08: d <= 8'h00; 15'h5F09: d <= 8'h00; 15'h5F0A: d <= 8'h00; 15'h5F0B: d <= 8'h00;
                15'h5F0C: d <= 8'h00; 15'h5F0D: d <= 8'h00; 15'h5F0E: d <= 8'h00; 15'h5F0F: d <= 8'h00;
                15'h5F10: d <= 8'h00; 15'h5F11: d <= 8'h00; 15'h5F12: d <= 8'h00; 15'h5F13: d <= 8'h00;
                15'h5F14: d <= 8'h00; 15'h5F15: d <= 8'h00; 15'h5F16: d <= 8'h00; 15'h5F17: d <= 8'h00;
                15'h5F18: d <= 8'h00; 15'h5F19: d <= 8'h00; 15'h5F1A: d <= 8'h00; 15'h5F1B: d <= 8'h00;
                15'h5F1C: d <= 8'h00; 15'h5F1D: d <= 8'h00; 15'h5F1E: d <= 8'h00; 15'h5F1F: d <= 8'h00;
                15'h5F20: d <= 8'h00; 15'h5F21: d <= 8'h00; 15'h5F22: d <= 8'h00; 15'h5F23: d <= 8'h00;
                15'h5F24: d <= 8'h00; 15'h5F25: d <= 8'h00; 15'h5F26: d <= 8'h00; 15'h5F27: d <= 8'h00;
                15'h5F28: d <= 8'h00; 15'h5F29: d <= 8'h00; 15'h5F2A: d <= 8'h00; 15'h5F2B: d <= 8'h00;
                15'h5F2C: d <= 8'h00; 15'h5F2D: d <= 8'h00; 15'h5F2E: d <= 8'h00; 15'h5F2F: d <= 8'h7B;
                15'h5F30: d <= 8'h00; 15'h5F31: d <= 8'h00; 15'h5F32: d <= 8'h00; 15'h5F33: d <= 8'h00;
                15'h5F34: d <= 8'h00; 15'h5F35: d <= 8'h00; 15'h5F36: d <= 8'h00; 15'h5F37: d <= 8'h00;
                15'h5F38: d <= 8'h00; 15'h5F39: d <= 8'h00; 15'h5F3A: d <= 8'h00; 15'h5F3B: d <= 8'h00;
                15'h5F3C: d <= 8'h00; 15'h5F3D: d <= 8'h00; 15'h5F3E: d <= 8'h00; 15'h5F3F: d <= 8'h00;
                15'h5F40: d <= 8'h00; 15'h5F41: d <= 8'h00; 15'h5F42: d <= 8'h00; 15'h5F43: d <= 8'h00;
                15'h5F44: d <= 8'h00; 15'h5F45: d <= 8'h00; 15'h5F46: d <= 8'h00; 15'h5F47: d <= 8'h00;
                15'h5F48: d <= 8'h00; 15'h5F49: d <= 8'h00; 15'h5F4A: d <= 8'h00; 15'h5F4B: d <= 8'h00;
                15'h5F4C: d <= 8'h00; 15'h5F4D: d <= 8'h00; 15'h5F4E: d <= 8'h00; 15'h5F4F: d <= 8'h00;
                15'h5F50: d <= 8'h00; 15'h5F51: d <= 8'h00; 15'h5F52: d <= 8'h00; 15'h5F53: d <= 8'h00;
                15'h5F54: d <= 8'h00; 15'h5F55: d <= 8'h00; 15'h5F56: d <= 8'h00; 15'h5F57: d <= 8'h00;
                15'h5F58: d <= 8'h45; 15'h5F59: d <= 8'h35; 15'h5F5A: d <= 8'h32; 15'h5F5B: d <= 8'h00;
                15'h5F5C: d <= 8'h00; 15'h5F5D: d <= 8'h00; 15'h5F5E: d <= 8'h00; 15'h5F5F: d <= 8'h00;
                15'h5F60: d <= 8'h00; 15'h5F61: d <= 8'h00; 15'h5F62: d <= 8'h00; 15'h5F63: d <= 8'h00;
                15'h5F64: d <= 8'h00; 15'h5F65: d <= 8'h00; 15'h5F66: d <= 8'h00; 15'h5F67: d <= 8'h00;
                15'h5F68: d <= 8'h00; 15'h5F69: d <= 8'h00; 15'h5F6A: d <= 8'h00; 15'h5F6B: d <= 8'h00;
                15'h5F6C: d <= 8'h00; 15'h5F6D: d <= 8'h00; 15'h5F6E: d <= 8'h00; 15'h5F6F: d <= 8'h00;
                15'h5F70: d <= 8'h00; 15'h5F71: d <= 8'h00; 15'h5F72: d <= 8'h00; 15'h5F73: d <= 8'h00;
                15'h5F74: d <= 8'h00; 15'h5F75: d <= 8'h00; 15'h5F76: d <= 8'h00; 15'h5F77: d <= 8'h00;
                15'h5F78: d <= 8'h00; 15'h5F79: d <= 8'h00; 15'h5F7A: d <= 8'h00; 15'h5F7B: d <= 8'h00;
                15'h5F7C: d <= 8'h00; 15'h5F7D: d <= 8'h00; 15'h5F7E: d <= 8'h00; 15'h5F7F: d <= 8'hE0;
                15'h5F80: d <= 8'h10; 15'h5F81: d <= 8'h15; 15'h5F82: d <= 8'h1A; 15'h5F83: d <= 8'h1F;
                15'h5F84: d <= 8'h20; 15'h5F85: d <= 8'h25; 15'h5F86: d <= 8'h2A; 15'h5F87: d <= 8'h2F;
                15'h5F88: d <= 8'h34; 15'h5F89: d <= 8'h38; 15'h5F8A: d <= 8'h3C; 15'h5F8B: d <= 8'h31;
                15'h5F8C: d <= 8'h39; 15'h5F8D: d <= 8'h3D; 15'h5F8E: d <= 8'h32; 15'h5F8F: d <= 8'h36;
                15'h5F90: d <= 8'h3E; 15'h5F91: d <= 8'h33; 15'h5F92: d <= 8'h37; 15'h5F93: d <= 8'h3B;
                15'h5F94: d <= 8'h44; 15'h5F95: d <= 8'h48; 15'h5F96: d <= 8'h4C; 15'h5F97: d <= 8'h41;
                15'h5F98: d <= 8'h49; 15'h5F99: d <= 8'h4D; 15'h5F9A: d <= 8'h42; 15'h5F9B: d <= 8'h46;
                15'h5F9C: d <= 8'h4E; 15'h5F9D: d <= 8'h43; 15'h5F9E: d <= 8'h47; 15'h5F9F: d <= 8'h4B;
                15'h5FA0: d <= 8'h50; 15'h5FA1: d <= 8'h55; 15'h5FA2: d <= 8'h5A; 15'h5FA3: d <= 8'h5F;
                15'h5FA4: d <= 8'h60; 15'h5FA5: d <= 8'h65; 15'h5FA6: d <= 8'h6A; 15'h5FA7: d <= 8'h6F;
                15'h5FA8: d <= 8'h74; 15'h5FA9: d <= 8'h78; 15'h5FAA: d <= 8'h7C; 15'h5FAB: d <= 8'h71;
                15'h5FAC: d <= 8'h79; 15'h5FAD: d <= 8'h7D; 15'h5FAE: d <= 8'h72; 15'h5FAF: d <= 8'h76;
                15'h5FB0: d <= 8'h7E; 15'h5FB1: d <= 8'h73; 15'h5FB2: d <= 8'h77; 15'h5FB3: d <= 8'h7B;
                15'h5FB4: d <= 8'h84; 15'h5FB5: d <= 8'h88; 15'h5FB6: d <= 8'h8C; 15'h5FB7: d <= 8'h81;
                15'h5FB8: d <= 8'h89; 15'h5FB9: d <= 8'h8D; 15'h5FBA: d <= 8'h82; 15'h5FBB: d <= 8'h86;
                15'h5FBC: d <= 8'h8E; 15'h5FBD: d <= 8'h83; 15'h5FBE: d <= 8'h87; 15'h5FBF: d <= 8'h8B;
                15'h5FC0: d <= 8'h90; 15'h5FC1: d <= 8'h95; 15'h5FC2: d <= 8'h9A; 15'h5FC3: d <= 8'h9F;
                15'h5FC4: d <= 8'hA4; 15'h5FC5: d <= 8'hA8; 15'h5FC6: d <= 8'hAC; 15'h5FC7: d <= 8'hA1;
                15'h5FC8: d <= 8'hA9; 15'h5FC9: d <= 8'hAD; 15'h5FCA: d <= 8'hA2; 15'h5FCB: d <= 8'hA6;
                15'h5FCC: d <= 8'hAE; 15'h5FCD: d <= 8'hA3; 15'h5FCE: d <= 8'hA7; 15'h5FCF: d <= 8'hAB;
                15'h5FD0: d <= 8'hB4; 15'h5FD1: d <= 8'hB8; 15'h5FD2: d <= 8'hBC; 15'h5FD3: d <= 8'hB1;
                15'h5FD4: d <= 8'hB9; 15'h5FD5: d <= 8'hBD; 15'h5FD6: d <= 8'hB2; 15'h5FD7: d <= 8'hB6;
                15'h5FD8: d <= 8'hBE; 15'h5FD9: d <= 8'hB3; 15'h5FDA: d <= 8'hB7; 15'h5FDB: d <= 8'hBB;
                15'h5FDC: d <= 8'hC4; 15'h5FDD: d <= 8'hC8; 15'h5FDE: d <= 8'hCC; 15'h5FDF: d <= 8'hC1;
                15'h5FE0: d <= 8'hC9; 15'h5FE1: d <= 8'hCD; 15'h5FE2: d <= 8'hC2; 15'h5FE3: d <= 8'hC6;
                15'h5FE4: d <= 8'hCE; 15'h5FE5: d <= 8'hC3; 15'h5FE6: d <= 8'hC7; 15'h5FE7: d <= 8'hCB;
                15'h5FE8: d <= 8'hC0; 15'h5FE9: d <= 8'hC5; 15'h5FEA: d <= 8'hCA; 15'h5FEB: d <= 8'hCF;
                15'h5FEC: d <= 8'hD0; 15'h5FED: d <= 8'hD5; 15'h5FEE: d <= 8'hDA; 15'h5FEF: d <= 8'hDF;
                15'h5FF0: d <= 8'h74; 15'h5FF1: d <= 8'h78; 15'h5FF2: d <= 8'h7C; 15'h5FF3: d <= 8'h71;
                15'h5FF4: d <= 8'h79; 15'h5FF5: d <= 8'h7D; 15'h5FF6: d <= 8'h72; 15'h5FF7: d <= 8'h76;
                15'h5FF8: d <= 8'h7E; 15'h5FF9: d <= 8'h73; 15'h5FFA: d <= 8'h77; 15'h5FFB: d <= 8'h7B;
                15'h5FFC: d <= 8'hA0; 15'h5FFD: d <= 8'hA5; 15'h5FFE: d <= 8'hAA; 15'h5FFF: d <= 8'hAF;
                15'h6000: d <= 8'h00; 15'h6001: d <= 8'h00; 15'h6002: d <= 8'h00; 15'h6003: d <= 8'h00;
                15'h6004: d <= 8'h00; 15'h6005: d <= 8'h00; 15'h6006: d <= 8'h00; 15'h6007: d <= 8'h00;
                15'h6008: d <= 8'h00; 15'h6009: d <= 8'h00; 15'h600A: d <= 8'h00; 15'h600B: d <= 8'h00;
                15'h600C: d <= 8'h00; 15'h600D: d <= 8'h00; 15'h600E: d <= 8'h00; 15'h600F: d <= 8'h00;
                15'h6010: d <= 8'h00; 15'h6011: d <= 8'h00; 15'h6012: d <= 8'h00; 15'h6013: d <= 8'h00;
                15'h6014: d <= 8'h00; 15'h6015: d <= 8'h00; 15'h6016: d <= 8'h00; 15'h6017: d <= 8'h00;
                15'h6018: d <= 8'h00; 15'h6019: d <= 8'h00; 15'h601A: d <= 8'h00; 15'h601B: d <= 8'h00;
                15'h601C: d <= 8'h00; 15'h601D: d <= 8'h00; 15'h601E: d <= 8'h00; 15'h601F: d <= 8'h00;
                15'h6020: d <= 8'h00; 15'h6021: d <= 8'h00; 15'h6022: d <= 8'h00; 15'h6023: d <= 8'h00;
                15'h6024: d <= 8'h00; 15'h6025: d <= 8'h00; 15'h6026: d <= 8'h00; 15'h6027: d <= 8'h00;
                15'h6028: d <= 8'h00; 15'h6029: d <= 8'h00; 15'h602A: d <= 8'h00; 15'h602B: d <= 8'h00;
                15'h602C: d <= 8'h00; 15'h602D: d <= 8'h00; 15'h602E: d <= 8'h00; 15'h602F: d <= 8'hAF;
                15'h6030: d <= 8'h00; 15'h6031: d <= 8'h00; 15'h6032: d <= 8'h00; 15'h6033: d <= 8'h00;
                15'h6034: d <= 8'h00; 15'h6035: d <= 8'h00; 15'h6036: d <= 8'h00; 15'h6037: d <= 8'h00;
                15'h6038: d <= 8'h00; 15'h6039: d <= 8'h00; 15'h603A: d <= 8'h00; 15'h603B: d <= 8'h00;
                15'h603C: d <= 8'h00; 15'h603D: d <= 8'h00; 15'h603E: d <= 8'h00; 15'h603F: d <= 8'h00;
                15'h6040: d <= 8'h00; 15'h6041: d <= 8'h00; 15'h6042: d <= 8'h00; 15'h6043: d <= 8'h00;
                15'h6044: d <= 8'h00; 15'h6045: d <= 8'h00; 15'h6046: d <= 8'h00; 15'h6047: d <= 8'h00;
                15'h6048: d <= 8'h00; 15'h6049: d <= 8'h00; 15'h604A: d <= 8'h00; 15'h604B: d <= 8'h00;
                15'h604C: d <= 8'h00; 15'h604D: d <= 8'h00; 15'h604E: d <= 8'h00; 15'h604F: d <= 8'h00;
                15'h6050: d <= 8'h00; 15'h6051: d <= 8'h00; 15'h6052: d <= 8'h00; 15'h6053: d <= 8'h00;
                15'h6054: d <= 8'h00; 15'h6055: d <= 8'h00; 15'h6056: d <= 8'h00; 15'h6057: d <= 8'h00;
                15'h6058: d <= 8'h45; 15'h6059: d <= 8'h35; 15'h605A: d <= 8'hAA; 15'h605B: d <= 8'h00;
                15'h605C: d <= 8'h00; 15'h605D: d <= 8'h00; 15'h605E: d <= 8'h00; 15'h605F: d <= 8'h00;
                15'h6060: d <= 8'h00; 15'h6061: d <= 8'h00; 15'h6062: d <= 8'h00; 15'h6063: d <= 8'h00;
                15'h6064: d <= 8'h00; 15'h6065: d <= 8'h00; 15'h6066: d <= 8'h00; 15'h6067: d <= 8'h00;
                15'h6068: d <= 8'h00; 15'h6069: d <= 8'h00; 15'h606A: d <= 8'h00; 15'h606B: d <= 8'h00;
                15'h606C: d <= 8'h00; 15'h606D: d <= 8'h00; 15'h606E: d <= 8'h00; 15'h606F: d <= 8'h00;
                15'h6070: d <= 8'h00; 15'h6071: d <= 8'h00; 15'h6072: d <= 8'h00; 15'h6073: d <= 8'h00;
                15'h6074: d <= 8'h00; 15'h6075: d <= 8'h00; 15'h6076: d <= 8'h00; 15'h6077: d <= 8'h00;
                15'h6078: d <= 8'h00; 15'h6079: d <= 8'h00; 15'h607A: d <= 8'h00; 15'h607B: d <= 8'h00;
                15'h607C: d <= 8'h00; 15'h607D: d <= 8'h00; 15'h607E: d <= 8'h00; 15'h607F: d <= 8'hE0;
                15'h6080: d <= 8'h10; 15'h6081: d <= 8'h15; 15'h6082: d <= 8'h1A; 15'h6083: d <= 8'h1F;
                15'h6084: d <= 8'h20; 15'h6085: d <= 8'h25; 15'h6086: d <= 8'h2A; 15'h6087: d <= 8'h2F;
                15'h6088: d <= 8'h34; 15'h6089: d <= 8'h38; 15'h608A: d <= 8'h3C; 15'h608B: d <= 8'h31;
                15'h608C: d <= 8'h39; 15'h608D: d <= 8'h3D; 15'h608E: d <= 8'h32; 15'h608F: d <= 8'h36;
                15'h6090: d <= 8'h3E; 15'h6091: d <= 8'h33; 15'h6092: d <= 8'h37; 15'h6093: d <= 8'h3B;
                15'h6094: d <= 8'h44; 15'h6095: d <= 8'h48; 15'h6096: d <= 8'h4C; 15'h6097: d <= 8'h41;
                15'h6098: d <= 8'h49; 15'h6099: d <= 8'h4D; 15'h609A: d <= 8'h42; 15'h609B: d <= 8'h46;
                15'h609C: d <= 8'h4E; 15'h609D: d <= 8'h43; 15'h609E: d <= 8'h47; 15'h609F: d <= 8'h4B;
                15'h60A0: d <= 8'h50; 15'h60A1: d <= 8'h55; 15'h60A2: d <= 8'h5A; 15'h60A3: d <= 8'h5F;
                15'h60A4: d <= 8'h60; 15'h60A5: d <= 8'h65; 15'h60A6: d <= 8'h6A; 15'h60A7: d <= 8'h6F;
                15'h60A8: d <= 8'h74; 15'h60A9: d <= 8'h78; 15'h60AA: d <= 8'h7C; 15'h60AB: d <= 8'h71;
                15'h60AC: d <= 8'h79; 15'h60AD: d <= 8'h7D; 15'h60AE: d <= 8'h72; 15'h60AF: d <= 8'h76;
                15'h60B0: d <= 8'h7E; 15'h60B1: d <= 8'h73; 15'h60B2: d <= 8'h77; 15'h60B3: d <= 8'h7B;
                15'h60B4: d <= 8'h84; 15'h60B5: d <= 8'h88; 15'h60B6: d <= 8'h8C; 15'h60B7: d <= 8'h81;
                15'h60B8: d <= 8'h89; 15'h60B9: d <= 8'h8D; 15'h60BA: d <= 8'h82; 15'h60BB: d <= 8'h86;
                15'h60BC: d <= 8'h8E; 15'h60BD: d <= 8'h83; 15'h60BE: d <= 8'h87; 15'h60BF: d <= 8'h8B;
                15'h60C0: d <= 8'h90; 15'h60C1: d <= 8'h95; 15'h60C2: d <= 8'h9A; 15'h60C3: d <= 8'h9F;
                15'h60C4: d <= 8'hA4; 15'h60C5: d <= 8'hA8; 15'h60C6: d <= 8'hAC; 15'h60C7: d <= 8'hA1;
                15'h60C8: d <= 8'hA9; 15'h60C9: d <= 8'hAD; 15'h60CA: d <= 8'hA2; 15'h60CB: d <= 8'hA6;
                15'h60CC: d <= 8'hAE; 15'h60CD: d <= 8'hA3; 15'h60CE: d <= 8'hA7; 15'h60CF: d <= 8'hAB;
                15'h60D0: d <= 8'hB4; 15'h60D1: d <= 8'hB8; 15'h60D2: d <= 8'hBC; 15'h60D3: d <= 8'hB1;
                15'h60D4: d <= 8'hB9; 15'h60D5: d <= 8'hBD; 15'h60D6: d <= 8'hB2; 15'h60D7: d <= 8'hB6;
                15'h60D8: d <= 8'hBE; 15'h60D9: d <= 8'hB3; 15'h60DA: d <= 8'hB7; 15'h60DB: d <= 8'hBB;
                15'h60DC: d <= 8'hC4; 15'h60DD: d <= 8'hC8; 15'h60DE: d <= 8'hCC; 15'h60DF: d <= 8'hC1;
                15'h60E0: d <= 8'hC9; 15'h60E1: d <= 8'hCD; 15'h60E2: d <= 8'hC2; 15'h60E3: d <= 8'hC6;
                15'h60E4: d <= 8'hCE; 15'h60E5: d <= 8'hC3; 15'h60E6: d <= 8'hC7; 15'h60E7: d <= 8'hCB;
                15'h60E8: d <= 8'hC0; 15'h60E9: d <= 8'hC5; 15'h60EA: d <= 8'hCA; 15'h60EB: d <= 8'hCF;
                15'h60EC: d <= 8'hD0; 15'h60ED: d <= 8'hD5; 15'h60EE: d <= 8'hDA; 15'h60EF: d <= 8'hDF;
                15'h60F0: d <= 8'h74; 15'h60F1: d <= 8'h78; 15'h60F2: d <= 8'h7C; 15'h60F3: d <= 8'h71;
                15'h60F4: d <= 8'h79; 15'h60F5: d <= 8'h7D; 15'h60F6: d <= 8'h72; 15'h60F7: d <= 8'h76;
                15'h60F8: d <= 8'h7E; 15'h60F9: d <= 8'h73; 15'h60FA: d <= 8'h77; 15'h60FB: d <= 8'h7B;
                15'h60FC: d <= 8'hA0; 15'h60FD: d <= 8'hA5; 15'h60FE: d <= 8'hAA; 15'h60FF: d <= 8'hAF;
                15'h6100: d <= 8'h00; 15'h6101: d <= 8'h00; 15'h6102: d <= 8'h00; 15'h6103: d <= 8'h00;
                15'h6104: d <= 8'h00; 15'h6105: d <= 8'h00; 15'h6106: d <= 8'h00; 15'h6107: d <= 8'h00;
                15'h6108: d <= 8'h00; 15'h6109: d <= 8'h00; 15'h610A: d <= 8'h00; 15'h610B: d <= 8'h00;
                15'h610C: d <= 8'h00; 15'h610D: d <= 8'h00; 15'h610E: d <= 8'h00; 15'h610F: d <= 8'h00;
                15'h6110: d <= 8'h00; 15'h6111: d <= 8'h00; 15'h6112: d <= 8'h00; 15'h6113: d <= 8'h00;
                15'h6114: d <= 8'h00; 15'h6115: d <= 8'h00; 15'h6116: d <= 8'h00; 15'h6117: d <= 8'h00;
                15'h6118: d <= 8'h00; 15'h6119: d <= 8'h00; 15'h611A: d <= 8'h00; 15'h611B: d <= 8'h00;
                15'h611C: d <= 8'h00; 15'h611D: d <= 8'h00; 15'h611E: d <= 8'h00; 15'h611F: d <= 8'h00;
                15'h6120: d <= 8'h00; 15'h6121: d <= 8'h00; 15'h6122: d <= 8'h00; 15'h6123: d <= 8'h00;
                15'h6124: d <= 8'h00; 15'h6125: d <= 8'h00; 15'h6126: d <= 8'h00; 15'h6127: d <= 8'h00;
                15'h6128: d <= 8'h00; 15'h6129: d <= 8'h00; 15'h612A: d <= 8'h00; 15'h612B: d <= 8'h00;
                15'h612C: d <= 8'h00; 15'h612D: d <= 8'h00; 15'h612E: d <= 8'h00; 15'h612F: d <= 8'hAF;
                15'h6130: d <= 8'h00; 15'h6131: d <= 8'h00; 15'h6132: d <= 8'h00; 15'h6133: d <= 8'h00;
                15'h6134: d <= 8'h00; 15'h6135: d <= 8'h00; 15'h6136: d <= 8'h00; 15'h6137: d <= 8'h00;
                15'h6138: d <= 8'h00; 15'h6139: d <= 8'h00; 15'h613A: d <= 8'h00; 15'h613B: d <= 8'h00;
                15'h613C: d <= 8'h00; 15'h613D: d <= 8'h00; 15'h613E: d <= 8'h00; 15'h613F: d <= 8'h00;
                15'h6140: d <= 8'h00; 15'h6141: d <= 8'h00; 15'h6142: d <= 8'h00; 15'h6143: d <= 8'h00;
                15'h6144: d <= 8'h00; 15'h6145: d <= 8'h00; 15'h6146: d <= 8'h00; 15'h6147: d <= 8'h00;
                15'h6148: d <= 8'h00; 15'h6149: d <= 8'h00; 15'h614A: d <= 8'h00; 15'h614B: d <= 8'h00;
                15'h614C: d <= 8'h00; 15'h614D: d <= 8'h00; 15'h614E: d <= 8'h00; 15'h614F: d <= 8'h00;
                15'h6150: d <= 8'h00; 15'h6151: d <= 8'h00; 15'h6152: d <= 8'h00; 15'h6153: d <= 8'h00;
                15'h6154: d <= 8'h00; 15'h6155: d <= 8'h00; 15'h6156: d <= 8'h00; 15'h6157: d <= 8'h00;
                15'h6158: d <= 8'h45; 15'h6159: d <= 8'h35; 15'h615A: d <= 8'hAA; 15'h615B: d <= 8'h00;
                15'h615C: d <= 8'h00; 15'h615D: d <= 8'h00; 15'h615E: d <= 8'h00; 15'h615F: d <= 8'h00;
                15'h6160: d <= 8'h00; 15'h6161: d <= 8'h00; 15'h6162: d <= 8'h00; 15'h6163: d <= 8'h00;
                15'h6164: d <= 8'h00; 15'h6165: d <= 8'h00; 15'h6166: d <= 8'h00; 15'h6167: d <= 8'h00;
                15'h6168: d <= 8'h00; 15'h6169: d <= 8'h00; 15'h616A: d <= 8'h00; 15'h616B: d <= 8'h00;
                15'h616C: d <= 8'h00; 15'h616D: d <= 8'h00; 15'h616E: d <= 8'h00; 15'h616F: d <= 8'h00;
                15'h6170: d <= 8'h00; 15'h6171: d <= 8'h00; 15'h6172: d <= 8'h00; 15'h6173: d <= 8'h00;
                15'h6174: d <= 8'h00; 15'h6175: d <= 8'h00; 15'h6176: d <= 8'h00; 15'h6177: d <= 8'h00;
                15'h6178: d <= 8'h00; 15'h6179: d <= 8'h00; 15'h617A: d <= 8'h00; 15'h617B: d <= 8'h00;
                15'h617C: d <= 8'h00; 15'h617D: d <= 8'h00; 15'h617E: d <= 8'h00; 15'h617F: d <= 8'hE0;
                15'h6180: d <= 8'h10; 15'h6181: d <= 8'h15; 15'h6182: d <= 8'h1A; 15'h6183: d <= 8'h1F;
                15'h6184: d <= 8'h20; 15'h6185: d <= 8'h25; 15'h6186: d <= 8'h2A; 15'h6187: d <= 8'h2F;
                15'h6188: d <= 8'h34; 15'h6189: d <= 8'h38; 15'h618A: d <= 8'h3C; 15'h618B: d <= 8'h31;
                15'h618C: d <= 8'h39; 15'h618D: d <= 8'h3D; 15'h618E: d <= 8'h32; 15'h618F: d <= 8'h36;
                15'h6190: d <= 8'h3E; 15'h6191: d <= 8'h33; 15'h6192: d <= 8'h37; 15'h6193: d <= 8'h3B;
                15'h6194: d <= 8'h44; 15'h6195: d <= 8'h48; 15'h6196: d <= 8'h4C; 15'h6197: d <= 8'h41;
                15'h6198: d <= 8'h49; 15'h6199: d <= 8'h4D; 15'h619A: d <= 8'h42; 15'h619B: d <= 8'h46;
                15'h619C: d <= 8'h4E; 15'h619D: d <= 8'h43; 15'h619E: d <= 8'h47; 15'h619F: d <= 8'h4B;
                15'h61A0: d <= 8'h50; 15'h61A1: d <= 8'h55; 15'h61A2: d <= 8'h5A; 15'h61A3: d <= 8'h5F;
                15'h61A4: d <= 8'h60; 15'h61A5: d <= 8'h65; 15'h61A6: d <= 8'h6A; 15'h61A7: d <= 8'h6F;
                15'h61A8: d <= 8'h74; 15'h61A9: d <= 8'h78; 15'h61AA: d <= 8'h7C; 15'h61AB: d <= 8'h71;
                15'h61AC: d <= 8'h79; 15'h61AD: d <= 8'h7D; 15'h61AE: d <= 8'h72; 15'h61AF: d <= 8'h76;
                15'h61B0: d <= 8'h7E; 15'h61B1: d <= 8'h73; 15'h61B2: d <= 8'h77; 15'h61B3: d <= 8'h7B;
                15'h61B4: d <= 8'h84; 15'h61B5: d <= 8'h88; 15'h61B6: d <= 8'h8C; 15'h61B7: d <= 8'h81;
                15'h61B8: d <= 8'h89; 15'h61B9: d <= 8'h8D; 15'h61BA: d <= 8'h82; 15'h61BB: d <= 8'h86;
                15'h61BC: d <= 8'h8E; 15'h61BD: d <= 8'h83; 15'h61BE: d <= 8'h87; 15'h61BF: d <= 8'h8B;
                15'h61C0: d <= 8'h90; 15'h61C1: d <= 8'h95; 15'h61C2: d <= 8'h9A; 15'h61C3: d <= 8'h9F;
                15'h61C4: d <= 8'hA4; 15'h61C5: d <= 8'hA8; 15'h61C6: d <= 8'hAC; 15'h61C7: d <= 8'hA1;
                15'h61C8: d <= 8'hA9; 15'h61C9: d <= 8'hAD; 15'h61CA: d <= 8'hA2; 15'h61CB: d <= 8'hA6;
                15'h61CC: d <= 8'hAE; 15'h61CD: d <= 8'hA3; 15'h61CE: d <= 8'hA7; 15'h61CF: d <= 8'hAB;
                15'h61D0: d <= 8'hB4; 15'h61D1: d <= 8'hB8; 15'h61D2: d <= 8'hBC; 15'h61D3: d <= 8'hB1;
                15'h61D4: d <= 8'hB9; 15'h61D5: d <= 8'hBD; 15'h61D6: d <= 8'hB2; 15'h61D7: d <= 8'hB6;
                15'h61D8: d <= 8'hBE; 15'h61D9: d <= 8'hB3; 15'h61DA: d <= 8'hB7; 15'h61DB: d <= 8'hBB;
                15'h61DC: d <= 8'hC4; 15'h61DD: d <= 8'hC8; 15'h61DE: d <= 8'hCC; 15'h61DF: d <= 8'hC1;
                15'h61E0: d <= 8'hC9; 15'h61E1: d <= 8'hCD; 15'h61E2: d <= 8'hC2; 15'h61E3: d <= 8'hC6;
                15'h61E4: d <= 8'hCE; 15'h61E5: d <= 8'hC3; 15'h61E6: d <= 8'hC7; 15'h61E7: d <= 8'hCB;
                15'h61E8: d <= 8'hC0; 15'h61E9: d <= 8'hC5; 15'h61EA: d <= 8'hCA; 15'h61EB: d <= 8'hCF;
                15'h61EC: d <= 8'hD0; 15'h61ED: d <= 8'hD5; 15'h61EE: d <= 8'hDA; 15'h61EF: d <= 8'hDF;
                15'h61F0: d <= 8'h74; 15'h61F1: d <= 8'h78; 15'h61F2: d <= 8'h7C; 15'h61F3: d <= 8'h71;
                15'h61F4: d <= 8'h79; 15'h61F5: d <= 8'h7D; 15'h61F6: d <= 8'h72; 15'h61F7: d <= 8'h76;
                15'h61F8: d <= 8'h7E; 15'h61F9: d <= 8'h73; 15'h61FA: d <= 8'h77; 15'h61FB: d <= 8'h7B;
                15'h61FC: d <= 8'hA0; 15'h61FD: d <= 8'hA5; 15'h61FE: d <= 8'hAA; 15'h61FF: d <= 8'hAF;
                15'h6200: d <= 8'h00; 15'h6201: d <= 8'h00; 15'h6202: d <= 8'h00; 15'h6203: d <= 8'h00;
                15'h6204: d <= 8'h00; 15'h6205: d <= 8'h00; 15'h6206: d <= 8'h00; 15'h6207: d <= 8'h00;
                15'h6208: d <= 8'h00; 15'h6209: d <= 8'h00; 15'h620A: d <= 8'h00; 15'h620B: d <= 8'h00;
                15'h620C: d <= 8'h00; 15'h620D: d <= 8'h00; 15'h620E: d <= 8'h00; 15'h620F: d <= 8'h00;
                15'h6210: d <= 8'h00; 15'h6211: d <= 8'h00; 15'h6212: d <= 8'h00; 15'h6213: d <= 8'h00;
                15'h6214: d <= 8'h00; 15'h6215: d <= 8'h00; 15'h6216: d <= 8'h00; 15'h6217: d <= 8'h00;
                15'h6218: d <= 8'h00; 15'h6219: d <= 8'h00; 15'h621A: d <= 8'h00; 15'h621B: d <= 8'h00;
                15'h621C: d <= 8'h00; 15'h621D: d <= 8'h00; 15'h621E: d <= 8'h00; 15'h621F: d <= 8'h00;
                15'h6220: d <= 8'h00; 15'h6221: d <= 8'h00; 15'h6222: d <= 8'h00; 15'h6223: d <= 8'h00;
                15'h6224: d <= 8'h00; 15'h6225: d <= 8'h00; 15'h6226: d <= 8'h00; 15'h6227: d <= 8'h00;
                15'h6228: d <= 8'h00; 15'h6229: d <= 8'h00; 15'h622A: d <= 8'h00; 15'h622B: d <= 8'h00;
                15'h622C: d <= 8'h00; 15'h622D: d <= 8'h00; 15'h622E: d <= 8'h00; 15'h622F: d <= 8'hAF;
                15'h6230: d <= 8'h00; 15'h6231: d <= 8'h00; 15'h6232: d <= 8'h00; 15'h6233: d <= 8'h00;
                15'h6234: d <= 8'h00; 15'h6235: d <= 8'h00; 15'h6236: d <= 8'h00; 15'h6237: d <= 8'h00;
                15'h6238: d <= 8'h00; 15'h6239: d <= 8'h00; 15'h623A: d <= 8'h00; 15'h623B: d <= 8'h00;
                15'h623C: d <= 8'h00; 15'h623D: d <= 8'h00; 15'h623E: d <= 8'h00; 15'h623F: d <= 8'h00;
                15'h6240: d <= 8'h00; 15'h6241: d <= 8'h00; 15'h6242: d <= 8'h00; 15'h6243: d <= 8'h00;
                15'h6244: d <= 8'h00; 15'h6245: d <= 8'h00; 15'h6246: d <= 8'h00; 15'h6247: d <= 8'h00;
                15'h6248: d <= 8'h00; 15'h6249: d <= 8'h00; 15'h624A: d <= 8'h00; 15'h624B: d <= 8'h00;
                15'h624C: d <= 8'h00; 15'h624D: d <= 8'h00; 15'h624E: d <= 8'h00; 15'h624F: d <= 8'h00;
                15'h6250: d <= 8'h00; 15'h6251: d <= 8'h00; 15'h6252: d <= 8'h00; 15'h6253: d <= 8'h00;
                15'h6254: d <= 8'h00; 15'h6255: d <= 8'h00; 15'h6256: d <= 8'h00; 15'h6257: d <= 8'h00;
                15'h6258: d <= 8'h45; 15'h6259: d <= 8'h35; 15'h625A: d <= 8'hAA; 15'h625B: d <= 8'h00;
                15'h625C: d <= 8'h00; 15'h625D: d <= 8'h00; 15'h625E: d <= 8'h00; 15'h625F: d <= 8'h00;
                15'h6260: d <= 8'h00; 15'h6261: d <= 8'h00; 15'h6262: d <= 8'h00; 15'h6263: d <= 8'h00;
                15'h6264: d <= 8'h00; 15'h6265: d <= 8'h00; 15'h6266: d <= 8'h00; 15'h6267: d <= 8'h00;
                15'h6268: d <= 8'h00; 15'h6269: d <= 8'h00; 15'h626A: d <= 8'h00; 15'h626B: d <= 8'h00;
                15'h626C: d <= 8'h00; 15'h626D: d <= 8'h00; 15'h626E: d <= 8'h00; 15'h626F: d <= 8'h00;
                15'h6270: d <= 8'h00; 15'h6271: d <= 8'h00; 15'h6272: d <= 8'h00; 15'h6273: d <= 8'h00;
                15'h6274: d <= 8'h00; 15'h6275: d <= 8'h00; 15'h6276: d <= 8'h00; 15'h6277: d <= 8'h00;
                15'h6278: d <= 8'h00; 15'h6279: d <= 8'h00; 15'h627A: d <= 8'h00; 15'h627B: d <= 8'h00;
                15'h627C: d <= 8'h00; 15'h627D: d <= 8'h00; 15'h627E: d <= 8'h00; 15'h627F: d <= 8'hE0;
                15'h6280: d <= 8'h10; 15'h6281: d <= 8'h15; 15'h6282: d <= 8'h1A; 15'h6283: d <= 8'h1F;
                15'h6284: d <= 8'h20; 15'h6285: d <= 8'h25; 15'h6286: d <= 8'h2A; 15'h6287: d <= 8'h2F;
                15'h6288: d <= 8'h34; 15'h6289: d <= 8'h38; 15'h628A: d <= 8'h3C; 15'h628B: d <= 8'h31;
                15'h628C: d <= 8'h39; 15'h628D: d <= 8'h3D; 15'h628E: d <= 8'h32; 15'h628F: d <= 8'h36;
                15'h6290: d <= 8'h3E; 15'h6291: d <= 8'h33; 15'h6292: d <= 8'h37; 15'h6293: d <= 8'h3B;
                15'h6294: d <= 8'h44; 15'h6295: d <= 8'h48; 15'h6296: d <= 8'h4C; 15'h6297: d <= 8'h41;
                15'h6298: d <= 8'h49; 15'h6299: d <= 8'h4D; 15'h629A: d <= 8'h42; 15'h629B: d <= 8'h46;
                15'h629C: d <= 8'h4E; 15'h629D: d <= 8'h43; 15'h629E: d <= 8'h47; 15'h629F: d <= 8'h4B;
                15'h62A0: d <= 8'h50; 15'h62A1: d <= 8'h55; 15'h62A2: d <= 8'h5A; 15'h62A3: d <= 8'h5F;
                15'h62A4: d <= 8'h60; 15'h62A5: d <= 8'h65; 15'h62A6: d <= 8'h6A; 15'h62A7: d <= 8'h6F;
                15'h62A8: d <= 8'h74; 15'h62A9: d <= 8'h78; 15'h62AA: d <= 8'h7C; 15'h62AB: d <= 8'h71;
                15'h62AC: d <= 8'h79; 15'h62AD: d <= 8'h7D; 15'h62AE: d <= 8'h72; 15'h62AF: d <= 8'h76;
                15'h62B0: d <= 8'h7E; 15'h62B1: d <= 8'h73; 15'h62B2: d <= 8'h77; 15'h62B3: d <= 8'h7B;
                15'h62B4: d <= 8'h84; 15'h62B5: d <= 8'h88; 15'h62B6: d <= 8'h8C; 15'h62B7: d <= 8'h81;
                15'h62B8: d <= 8'h89; 15'h62B9: d <= 8'h8D; 15'h62BA: d <= 8'h82; 15'h62BB: d <= 8'h86;
                15'h62BC: d <= 8'h8E; 15'h62BD: d <= 8'h83; 15'h62BE: d <= 8'h87; 15'h62BF: d <= 8'h8B;
                15'h62C0: d <= 8'h90; 15'h62C1: d <= 8'h95; 15'h62C2: d <= 8'h9A; 15'h62C3: d <= 8'h9F;
                15'h62C4: d <= 8'hA4; 15'h62C5: d <= 8'hA8; 15'h62C6: d <= 8'hAC; 15'h62C7: d <= 8'hA1;
                15'h62C8: d <= 8'hA9; 15'h62C9: d <= 8'hAD; 15'h62CA: d <= 8'hA2; 15'h62CB: d <= 8'hA6;
                15'h62CC: d <= 8'hAE; 15'h62CD: d <= 8'hA3; 15'h62CE: d <= 8'hA7; 15'h62CF: d <= 8'hAB;
                15'h62D0: d <= 8'hB4; 15'h62D1: d <= 8'hB8; 15'h62D2: d <= 8'hBC; 15'h62D3: d <= 8'hB1;
                15'h62D4: d <= 8'hB9; 15'h62D5: d <= 8'hBD; 15'h62D6: d <= 8'hB2; 15'h62D7: d <= 8'hB6;
                15'h62D8: d <= 8'hBE; 15'h62D9: d <= 8'hB3; 15'h62DA: d <= 8'hB7; 15'h62DB: d <= 8'hBB;
                15'h62DC: d <= 8'hC4; 15'h62DD: d <= 8'hC8; 15'h62DE: d <= 8'hCC; 15'h62DF: d <= 8'hC1;
                15'h62E0: d <= 8'hC9; 15'h62E1: d <= 8'hCD; 15'h62E2: d <= 8'hC2; 15'h62E3: d <= 8'hC6;
                15'h62E4: d <= 8'hCE; 15'h62E5: d <= 8'hC3; 15'h62E6: d <= 8'hC7; 15'h62E7: d <= 8'hCB;
                15'h62E8: d <= 8'hC0; 15'h62E9: d <= 8'hC5; 15'h62EA: d <= 8'hCA; 15'h62EB: d <= 8'hCF;
                15'h62EC: d <= 8'hD0; 15'h62ED: d <= 8'hD5; 15'h62EE: d <= 8'hDA; 15'h62EF: d <= 8'hDF;
                15'h62F0: d <= 8'h74; 15'h62F1: d <= 8'h78; 15'h62F2: d <= 8'h7C; 15'h62F3: d <= 8'h71;
                15'h62F4: d <= 8'h79; 15'h62F5: d <= 8'h7D; 15'h62F6: d <= 8'h72; 15'h62F7: d <= 8'h76;
                15'h62F8: d <= 8'h7E; 15'h62F9: d <= 8'h73; 15'h62FA: d <= 8'h77; 15'h62FB: d <= 8'h7B;
                15'h62FC: d <= 8'hA0; 15'h62FD: d <= 8'hA5; 15'h62FE: d <= 8'hAA; 15'h62FF: d <= 8'hAF;
                15'h6300: d <= 8'h00; 15'h6301: d <= 8'h00; 15'h6302: d <= 8'h00; 15'h6303: d <= 8'h00;
                15'h6304: d <= 8'h00; 15'h6305: d <= 8'h00; 15'h6306: d <= 8'h00; 15'h6307: d <= 8'h00;
                15'h6308: d <= 8'h00; 15'h6309: d <= 8'h00; 15'h630A: d <= 8'h00; 15'h630B: d <= 8'h00;
                15'h630C: d <= 8'h00; 15'h630D: d <= 8'h00; 15'h630E: d <= 8'h00; 15'h630F: d <= 8'h00;
                15'h6310: d <= 8'h00; 15'h6311: d <= 8'h00; 15'h6312: d <= 8'h00; 15'h6313: d <= 8'h00;
                15'h6314: d <= 8'h00; 15'h6315: d <= 8'h00; 15'h6316: d <= 8'h00; 15'h6317: d <= 8'h00;
                15'h6318: d <= 8'h00; 15'h6319: d <= 8'h00; 15'h631A: d <= 8'h00; 15'h631B: d <= 8'h00;
                15'h631C: d <= 8'h00; 15'h631D: d <= 8'h00; 15'h631E: d <= 8'h00; 15'h631F: d <= 8'h00;
                15'h6320: d <= 8'h00; 15'h6321: d <= 8'h00; 15'h6322: d <= 8'h00; 15'h6323: d <= 8'h00;
                15'h6324: d <= 8'h00; 15'h6325: d <= 8'h00; 15'h6326: d <= 8'h00; 15'h6327: d <= 8'h00;
                15'h6328: d <= 8'h00; 15'h6329: d <= 8'h00; 15'h632A: d <= 8'h00; 15'h632B: d <= 8'h00;
                15'h632C: d <= 8'h00; 15'h632D: d <= 8'h00; 15'h632E: d <= 8'h00; 15'h632F: d <= 8'hAF;
                15'h6330: d <= 8'h00; 15'h6331: d <= 8'h00; 15'h6332: d <= 8'h00; 15'h6333: d <= 8'h00;
                15'h6334: d <= 8'h00; 15'h6335: d <= 8'h00; 15'h6336: d <= 8'h00; 15'h6337: d <= 8'h00;
                15'h6338: d <= 8'h00; 15'h6339: d <= 8'h00; 15'h633A: d <= 8'h00; 15'h633B: d <= 8'h00;
                15'h633C: d <= 8'h00; 15'h633D: d <= 8'h00; 15'h633E: d <= 8'h00; 15'h633F: d <= 8'h00;
                15'h6340: d <= 8'h00; 15'h6341: d <= 8'h00; 15'h6342: d <= 8'h00; 15'h6343: d <= 8'h00;
                15'h6344: d <= 8'h00; 15'h6345: d <= 8'h00; 15'h6346: d <= 8'h00; 15'h6347: d <= 8'h00;
                15'h6348: d <= 8'h00; 15'h6349: d <= 8'h00; 15'h634A: d <= 8'h00; 15'h634B: d <= 8'h00;
                15'h634C: d <= 8'h00; 15'h634D: d <= 8'h00; 15'h634E: d <= 8'h00; 15'h634F: d <= 8'h00;
                15'h6350: d <= 8'h00; 15'h6351: d <= 8'h00; 15'h6352: d <= 8'h00; 15'h6353: d <= 8'h00;
                15'h6354: d <= 8'h00; 15'h6355: d <= 8'h00; 15'h6356: d <= 8'h00; 15'h6357: d <= 8'h00;
                15'h6358: d <= 8'h45; 15'h6359: d <= 8'h35; 15'h635A: d <= 8'hAA; 15'h635B: d <= 8'h00;
                15'h635C: d <= 8'h00; 15'h635D: d <= 8'h00; 15'h635E: d <= 8'h00; 15'h635F: d <= 8'h00;
                15'h6360: d <= 8'h00; 15'h6361: d <= 8'h00; 15'h6362: d <= 8'h00; 15'h6363: d <= 8'h00;
                15'h6364: d <= 8'h00; 15'h6365: d <= 8'h00; 15'h6366: d <= 8'h00; 15'h6367: d <= 8'h00;
                15'h6368: d <= 8'h00; 15'h6369: d <= 8'h00; 15'h636A: d <= 8'h00; 15'h636B: d <= 8'h00;
                15'h636C: d <= 8'h00; 15'h636D: d <= 8'h00; 15'h636E: d <= 8'h00; 15'h636F: d <= 8'h00;
                15'h6370: d <= 8'h00; 15'h6371: d <= 8'h00; 15'h6372: d <= 8'h00; 15'h6373: d <= 8'h00;
                15'h6374: d <= 8'h00; 15'h6375: d <= 8'h00; 15'h6376: d <= 8'h00; 15'h6377: d <= 8'h00;
                15'h6378: d <= 8'h00; 15'h6379: d <= 8'h00; 15'h637A: d <= 8'h00; 15'h637B: d <= 8'h00;
                15'h637C: d <= 8'h00; 15'h637D: d <= 8'h00; 15'h637E: d <= 8'h00; 15'h637F: d <= 8'hE0;
                15'h6380: d <= 8'h10; 15'h6381: d <= 8'h15; 15'h6382: d <= 8'h1A; 15'h6383: d <= 8'h1F;
                15'h6384: d <= 8'h20; 15'h6385: d <= 8'h25; 15'h6386: d <= 8'h2A; 15'h6387: d <= 8'h2F;
                15'h6388: d <= 8'h34; 15'h6389: d <= 8'h38; 15'h638A: d <= 8'h3C; 15'h638B: d <= 8'h31;
                15'h638C: d <= 8'h39; 15'h638D: d <= 8'h3D; 15'h638E: d <= 8'h32; 15'h638F: d <= 8'h36;
                15'h6390: d <= 8'h3E; 15'h6391: d <= 8'h33; 15'h6392: d <= 8'h37; 15'h6393: d <= 8'h3B;
                15'h6394: d <= 8'h44; 15'h6395: d <= 8'h48; 15'h6396: d <= 8'h4C; 15'h6397: d <= 8'h41;
                15'h6398: d <= 8'h49; 15'h6399: d <= 8'h4D; 15'h639A: d <= 8'h42; 15'h639B: d <= 8'h46;
                15'h639C: d <= 8'h4E; 15'h639D: d <= 8'h43; 15'h639E: d <= 8'h47; 15'h639F: d <= 8'h4B;
                15'h63A0: d <= 8'h50; 15'h63A1: d <= 8'h55; 15'h63A2: d <= 8'h5A; 15'h63A3: d <= 8'h5F;
                15'h63A4: d <= 8'h60; 15'h63A5: d <= 8'h65; 15'h63A6: d <= 8'h6A; 15'h63A7: d <= 8'h6F;
                15'h63A8: d <= 8'h74; 15'h63A9: d <= 8'h78; 15'h63AA: d <= 8'h7C; 15'h63AB: d <= 8'h71;
                15'h63AC: d <= 8'h79; 15'h63AD: d <= 8'h7D; 15'h63AE: d <= 8'h72; 15'h63AF: d <= 8'h76;
                15'h63B0: d <= 8'h7E; 15'h63B1: d <= 8'h73; 15'h63B2: d <= 8'h77; 15'h63B3: d <= 8'h7B;
                15'h63B4: d <= 8'h84; 15'h63B5: d <= 8'h88; 15'h63B6: d <= 8'h8C; 15'h63B7: d <= 8'h81;
                15'h63B8: d <= 8'h89; 15'h63B9: d <= 8'h8D; 15'h63BA: d <= 8'h82; 15'h63BB: d <= 8'h86;
                15'h63BC: d <= 8'h8E; 15'h63BD: d <= 8'h83; 15'h63BE: d <= 8'h87; 15'h63BF: d <= 8'h8B;
                15'h63C0: d <= 8'h90; 15'h63C1: d <= 8'h95; 15'h63C2: d <= 8'h9A; 15'h63C3: d <= 8'h9F;
                15'h63C4: d <= 8'hA4; 15'h63C5: d <= 8'hA8; 15'h63C6: d <= 8'hAC; 15'h63C7: d <= 8'hA1;
                15'h63C8: d <= 8'hA9; 15'h63C9: d <= 8'hAD; 15'h63CA: d <= 8'hA2; 15'h63CB: d <= 8'hA6;
                15'h63CC: d <= 8'hAE; 15'h63CD: d <= 8'hA3; 15'h63CE: d <= 8'hA7; 15'h63CF: d <= 8'hAB;
                15'h63D0: d <= 8'hB4; 15'h63D1: d <= 8'hB8; 15'h63D2: d <= 8'hBC; 15'h63D3: d <= 8'hB1;
                15'h63D4: d <= 8'hB9; 15'h63D5: d <= 8'hBD; 15'h63D6: d <= 8'hB2; 15'h63D7: d <= 8'hB6;
                15'h63D8: d <= 8'hBE; 15'h63D9: d <= 8'hB3; 15'h63DA: d <= 8'hB7; 15'h63DB: d <= 8'hBB;
                15'h63DC: d <= 8'hC4; 15'h63DD: d <= 8'hC8; 15'h63DE: d <= 8'hCC; 15'h63DF: d <= 8'hC1;
                15'h63E0: d <= 8'hC9; 15'h63E1: d <= 8'hCD; 15'h63E2: d <= 8'hC2; 15'h63E3: d <= 8'hC6;
                15'h63E4: d <= 8'hCE; 15'h63E5: d <= 8'hC3; 15'h63E6: d <= 8'hC7; 15'h63E7: d <= 8'hCB;
                15'h63E8: d <= 8'hC0; 15'h63E9: d <= 8'hC5; 15'h63EA: d <= 8'hCA; 15'h63EB: d <= 8'hCF;
                15'h63EC: d <= 8'hD0; 15'h63ED: d <= 8'hD5; 15'h63EE: d <= 8'hDA; 15'h63EF: d <= 8'hDF;
                15'h63F0: d <= 8'h74; 15'h63F1: d <= 8'h78; 15'h63F2: d <= 8'h7C; 15'h63F3: d <= 8'h71;
                15'h63F4: d <= 8'h79; 15'h63F5: d <= 8'h7D; 15'h63F6: d <= 8'h72; 15'h63F7: d <= 8'h76;
                15'h63F8: d <= 8'h7E; 15'h63F9: d <= 8'h73; 15'h63FA: d <= 8'h77; 15'h63FB: d <= 8'h7B;
                15'h63FC: d <= 8'hA0; 15'h63FD: d <= 8'hA5; 15'h63FE: d <= 8'hAA; 15'h63FF: d <= 8'hAF;
                15'h6400: d <= 8'h00; 15'h6401: d <= 8'h00; 15'h6402: d <= 8'h00; 15'h6403: d <= 8'h00;
                15'h6404: d <= 8'h00; 15'h6405: d <= 8'h00; 15'h6406: d <= 8'h00; 15'h6407: d <= 8'h00;
                15'h6408: d <= 8'h00; 15'h6409: d <= 8'h00; 15'h640A: d <= 8'h00; 15'h640B: d <= 8'h00;
                15'h640C: d <= 8'h00; 15'h640D: d <= 8'h00; 15'h640E: d <= 8'h00; 15'h640F: d <= 8'h00;
                15'h6410: d <= 8'h00; 15'h6411: d <= 8'h00; 15'h6412: d <= 8'h00; 15'h6413: d <= 8'h00;
                15'h6414: d <= 8'h00; 15'h6415: d <= 8'h00; 15'h6416: d <= 8'h00; 15'h6417: d <= 8'h00;
                15'h6418: d <= 8'h00; 15'h6419: d <= 8'h00; 15'h641A: d <= 8'h00; 15'h641B: d <= 8'h00;
                15'h641C: d <= 8'h00; 15'h641D: d <= 8'h00; 15'h641E: d <= 8'h00; 15'h641F: d <= 8'h00;
                15'h6420: d <= 8'h00; 15'h6421: d <= 8'h00; 15'h6422: d <= 8'h00; 15'h6423: d <= 8'h00;
                15'h6424: d <= 8'h00; 15'h6425: d <= 8'h00; 15'h6426: d <= 8'h00; 15'h6427: d <= 8'h00;
                15'h6428: d <= 8'h00; 15'h6429: d <= 8'h00; 15'h642A: d <= 8'h00; 15'h642B: d <= 8'h00;
                15'h642C: d <= 8'h00; 15'h642D: d <= 8'h00; 15'h642E: d <= 8'h00; 15'h642F: d <= 8'hAF;
                15'h6430: d <= 8'h00; 15'h6431: d <= 8'h00; 15'h6432: d <= 8'h00; 15'h6433: d <= 8'h00;
                15'h6434: d <= 8'h00; 15'h6435: d <= 8'h00; 15'h6436: d <= 8'h00; 15'h6437: d <= 8'h00;
                15'h6438: d <= 8'h00; 15'h6439: d <= 8'h00; 15'h643A: d <= 8'h00; 15'h643B: d <= 8'h00;
                15'h643C: d <= 8'h00; 15'h643D: d <= 8'h00; 15'h643E: d <= 8'h00; 15'h643F: d <= 8'h00;
                15'h6440: d <= 8'h00; 15'h6441: d <= 8'h00; 15'h6442: d <= 8'h00; 15'h6443: d <= 8'h00;
                15'h6444: d <= 8'h00; 15'h6445: d <= 8'h00; 15'h6446: d <= 8'h00; 15'h6447: d <= 8'h00;
                15'h6448: d <= 8'h00; 15'h6449: d <= 8'h00; 15'h644A: d <= 8'h00; 15'h644B: d <= 8'h00;
                15'h644C: d <= 8'h00; 15'h644D: d <= 8'h00; 15'h644E: d <= 8'h00; 15'h644F: d <= 8'h00;
                15'h6450: d <= 8'h00; 15'h6451: d <= 8'h00; 15'h6452: d <= 8'h00; 15'h6453: d <= 8'h00;
                15'h6454: d <= 8'h00; 15'h6455: d <= 8'h00; 15'h6456: d <= 8'h00; 15'h6457: d <= 8'h00;
                15'h6458: d <= 8'h45; 15'h6459: d <= 8'h35; 15'h645A: d <= 8'hAA; 15'h645B: d <= 8'h00;
                15'h645C: d <= 8'h00; 15'h645D: d <= 8'h00; 15'h645E: d <= 8'h00; 15'h645F: d <= 8'h00;
                15'h6460: d <= 8'h00; 15'h6461: d <= 8'h00; 15'h6462: d <= 8'h00; 15'h6463: d <= 8'h00;
                15'h6464: d <= 8'h00; 15'h6465: d <= 8'h00; 15'h6466: d <= 8'h00; 15'h6467: d <= 8'h00;
                15'h6468: d <= 8'h00; 15'h6469: d <= 8'h00; 15'h646A: d <= 8'h00; 15'h646B: d <= 8'h00;
                15'h646C: d <= 8'h00; 15'h646D: d <= 8'h00; 15'h646E: d <= 8'h00; 15'h646F: d <= 8'h00;
                15'h6470: d <= 8'h00; 15'h6471: d <= 8'h00; 15'h6472: d <= 8'h00; 15'h6473: d <= 8'h00;
                15'h6474: d <= 8'h00; 15'h6475: d <= 8'h00; 15'h6476: d <= 8'h00; 15'h6477: d <= 8'h00;
                15'h6478: d <= 8'h00; 15'h6479: d <= 8'h00; 15'h647A: d <= 8'h00; 15'h647B: d <= 8'h00;
                15'h647C: d <= 8'h00; 15'h647D: d <= 8'h00; 15'h647E: d <= 8'h00; 15'h647F: d <= 8'hE0;
                15'h6480: d <= 8'h10; 15'h6481: d <= 8'h15; 15'h6482: d <= 8'h1A; 15'h6483: d <= 8'h1F;
                15'h6484: d <= 8'h20; 15'h6485: d <= 8'h25; 15'h6486: d <= 8'h2A; 15'h6487: d <= 8'h2F;
                15'h6488: d <= 8'h34; 15'h6489: d <= 8'h38; 15'h648A: d <= 8'h3C; 15'h648B: d <= 8'h31;
                15'h648C: d <= 8'h39; 15'h648D: d <= 8'h3D; 15'h648E: d <= 8'h32; 15'h648F: d <= 8'h36;
                15'h6490: d <= 8'h3E; 15'h6491: d <= 8'h33; 15'h6492: d <= 8'h37; 15'h6493: d <= 8'h3B;
                15'h6494: d <= 8'h44; 15'h6495: d <= 8'h48; 15'h6496: d <= 8'h4C; 15'h6497: d <= 8'h41;
                15'h6498: d <= 8'h49; 15'h6499: d <= 8'h4D; 15'h649A: d <= 8'h42; 15'h649B: d <= 8'h46;
                15'h649C: d <= 8'h4E; 15'h649D: d <= 8'h43; 15'h649E: d <= 8'h47; 15'h649F: d <= 8'h4B;
                15'h64A0: d <= 8'h50; 15'h64A1: d <= 8'h55; 15'h64A2: d <= 8'h5A; 15'h64A3: d <= 8'h5F;
                15'h64A4: d <= 8'h60; 15'h64A5: d <= 8'h65; 15'h64A6: d <= 8'h6A; 15'h64A7: d <= 8'h6F;
                15'h64A8: d <= 8'h74; 15'h64A9: d <= 8'h78; 15'h64AA: d <= 8'h7C; 15'h64AB: d <= 8'h71;
                15'h64AC: d <= 8'h79; 15'h64AD: d <= 8'h7D; 15'h64AE: d <= 8'h72; 15'h64AF: d <= 8'h76;
                15'h64B0: d <= 8'h7E; 15'h64B1: d <= 8'h73; 15'h64B2: d <= 8'h77; 15'h64B3: d <= 8'h7B;
                15'h64B4: d <= 8'h84; 15'h64B5: d <= 8'h88; 15'h64B6: d <= 8'h8C; 15'h64B7: d <= 8'h81;
                15'h64B8: d <= 8'h89; 15'h64B9: d <= 8'h8D; 15'h64BA: d <= 8'h82; 15'h64BB: d <= 8'h86;
                15'h64BC: d <= 8'h8E; 15'h64BD: d <= 8'h83; 15'h64BE: d <= 8'h87; 15'h64BF: d <= 8'h8B;
                15'h64C0: d <= 8'h90; 15'h64C1: d <= 8'h95; 15'h64C2: d <= 8'h9A; 15'h64C3: d <= 8'h9F;
                15'h64C4: d <= 8'hA4; 15'h64C5: d <= 8'hA8; 15'h64C6: d <= 8'hAC; 15'h64C7: d <= 8'hA1;
                15'h64C8: d <= 8'hA9; 15'h64C9: d <= 8'hAD; 15'h64CA: d <= 8'hA2; 15'h64CB: d <= 8'hA6;
                15'h64CC: d <= 8'hAE; 15'h64CD: d <= 8'hA3; 15'h64CE: d <= 8'hA7; 15'h64CF: d <= 8'hAB;
                15'h64D0: d <= 8'hB4; 15'h64D1: d <= 8'hB8; 15'h64D2: d <= 8'hBC; 15'h64D3: d <= 8'hB1;
                15'h64D4: d <= 8'hB9; 15'h64D5: d <= 8'hBD; 15'h64D6: d <= 8'hB2; 15'h64D7: d <= 8'hB6;
                15'h64D8: d <= 8'hBE; 15'h64D9: d <= 8'hB3; 15'h64DA: d <= 8'hB7; 15'h64DB: d <= 8'hBB;
                15'h64DC: d <= 8'hC4; 15'h64DD: d <= 8'hC8; 15'h64DE: d <= 8'hCC; 15'h64DF: d <= 8'hC1;
                15'h64E0: d <= 8'hC9; 15'h64E1: d <= 8'hCD; 15'h64E2: d <= 8'hC2; 15'h64E3: d <= 8'hC6;
                15'h64E4: d <= 8'hCE; 15'h64E5: d <= 8'hC3; 15'h64E6: d <= 8'hC7; 15'h64E7: d <= 8'hCB;
                15'h64E8: d <= 8'hC0; 15'h64E9: d <= 8'hC5; 15'h64EA: d <= 8'hCA; 15'h64EB: d <= 8'hCF;
                15'h64EC: d <= 8'hD0; 15'h64ED: d <= 8'hD5; 15'h64EE: d <= 8'hDA; 15'h64EF: d <= 8'hDF;
                15'h64F0: d <= 8'h74; 15'h64F1: d <= 8'h78; 15'h64F2: d <= 8'h7C; 15'h64F3: d <= 8'h71;
                15'h64F4: d <= 8'h79; 15'h64F5: d <= 8'h7D; 15'h64F6: d <= 8'h72; 15'h64F7: d <= 8'h76;
                15'h64F8: d <= 8'h7E; 15'h64F9: d <= 8'h73; 15'h64FA: d <= 8'h77; 15'h64FB: d <= 8'h7B;
                15'h64FC: d <= 8'hA0; 15'h64FD: d <= 8'hA5; 15'h64FE: d <= 8'hAA; 15'h64FF: d <= 8'hAF;
                15'h6500: d <= 8'h00; 15'h6501: d <= 8'h00; 15'h6502: d <= 8'h00; 15'h6503: d <= 8'h00;
                15'h6504: d <= 8'h00; 15'h6505: d <= 8'h00; 15'h6506: d <= 8'h00; 15'h6507: d <= 8'h00;
                15'h6508: d <= 8'h00; 15'h6509: d <= 8'h00; 15'h650A: d <= 8'h00; 15'h650B: d <= 8'h00;
                15'h650C: d <= 8'h00; 15'h650D: d <= 8'h00; 15'h650E: d <= 8'h00; 15'h650F: d <= 8'h00;
                15'h6510: d <= 8'h00; 15'h6511: d <= 8'h00; 15'h6512: d <= 8'h00; 15'h6513: d <= 8'h00;
                15'h6514: d <= 8'h00; 15'h6515: d <= 8'h00; 15'h6516: d <= 8'h00; 15'h6517: d <= 8'h00;
                15'h6518: d <= 8'h00; 15'h6519: d <= 8'h00; 15'h651A: d <= 8'h00; 15'h651B: d <= 8'h00;
                15'h651C: d <= 8'h00; 15'h651D: d <= 8'h00; 15'h651E: d <= 8'h00; 15'h651F: d <= 8'h00;
                15'h6520: d <= 8'h00; 15'h6521: d <= 8'h00; 15'h6522: d <= 8'h00; 15'h6523: d <= 8'h00;
                15'h6524: d <= 8'h00; 15'h6525: d <= 8'h00; 15'h6526: d <= 8'h00; 15'h6527: d <= 8'h00;
                15'h6528: d <= 8'h00; 15'h6529: d <= 8'h00; 15'h652A: d <= 8'h00; 15'h652B: d <= 8'h00;
                15'h652C: d <= 8'h00; 15'h652D: d <= 8'h00; 15'h652E: d <= 8'h00; 15'h652F: d <= 8'hAF;
                15'h6530: d <= 8'h00; 15'h6531: d <= 8'h00; 15'h6532: d <= 8'h00; 15'h6533: d <= 8'h00;
                15'h6534: d <= 8'h00; 15'h6535: d <= 8'h00; 15'h6536: d <= 8'h00; 15'h6537: d <= 8'h00;
                15'h6538: d <= 8'h00; 15'h6539: d <= 8'h00; 15'h653A: d <= 8'h00; 15'h653B: d <= 8'h00;
                15'h653C: d <= 8'h00; 15'h653D: d <= 8'h00; 15'h653E: d <= 8'h00; 15'h653F: d <= 8'h00;
                15'h6540: d <= 8'h00; 15'h6541: d <= 8'h00; 15'h6542: d <= 8'h00; 15'h6543: d <= 8'h00;
                15'h6544: d <= 8'h00; 15'h6545: d <= 8'h00; 15'h6546: d <= 8'h00; 15'h6547: d <= 8'h00;
                15'h6548: d <= 8'h00; 15'h6549: d <= 8'h00; 15'h654A: d <= 8'h00; 15'h654B: d <= 8'h00;
                15'h654C: d <= 8'h00; 15'h654D: d <= 8'h00; 15'h654E: d <= 8'h00; 15'h654F: d <= 8'h00;
                15'h6550: d <= 8'h00; 15'h6551: d <= 8'h00; 15'h6552: d <= 8'h00; 15'h6553: d <= 8'h00;
                15'h6554: d <= 8'h00; 15'h6555: d <= 8'h00; 15'h6556: d <= 8'h00; 15'h6557: d <= 8'h00;
                15'h6558: d <= 8'h45; 15'h6559: d <= 8'h35; 15'h655A: d <= 8'hAA; 15'h655B: d <= 8'h00;
                15'h655C: d <= 8'h00; 15'h655D: d <= 8'h00; 15'h655E: d <= 8'h00; 15'h655F: d <= 8'h00;
                15'h6560: d <= 8'h00; 15'h6561: d <= 8'h00; 15'h6562: d <= 8'h00; 15'h6563: d <= 8'h00;
                15'h6564: d <= 8'h00; 15'h6565: d <= 8'h00; 15'h6566: d <= 8'h00; 15'h6567: d <= 8'h00;
                15'h6568: d <= 8'h00; 15'h6569: d <= 8'h00; 15'h656A: d <= 8'h00; 15'h656B: d <= 8'h00;
                15'h656C: d <= 8'h00; 15'h656D: d <= 8'h00; 15'h656E: d <= 8'h00; 15'h656F: d <= 8'h00;
                15'h6570: d <= 8'h00; 15'h6571: d <= 8'h00; 15'h6572: d <= 8'h00; 15'h6573: d <= 8'h00;
                15'h6574: d <= 8'h00; 15'h6575: d <= 8'h00; 15'h6576: d <= 8'h00; 15'h6577: d <= 8'h00;
                15'h6578: d <= 8'h00; 15'h6579: d <= 8'h00; 15'h657A: d <= 8'h00; 15'h657B: d <= 8'h00;
                15'h657C: d <= 8'h00; 15'h657D: d <= 8'h00; 15'h657E: d <= 8'h00; 15'h657F: d <= 8'hE0;
                15'h6580: d <= 8'h10; 15'h6581: d <= 8'h15; 15'h6582: d <= 8'h1A; 15'h6583: d <= 8'h1F;
                15'h6584: d <= 8'h20; 15'h6585: d <= 8'h25; 15'h6586: d <= 8'h2A; 15'h6587: d <= 8'h2F;
                15'h6588: d <= 8'h34; 15'h6589: d <= 8'h38; 15'h658A: d <= 8'h3C; 15'h658B: d <= 8'h31;
                15'h658C: d <= 8'h39; 15'h658D: d <= 8'h3D; 15'h658E: d <= 8'h32; 15'h658F: d <= 8'h36;
                15'h6590: d <= 8'h3E; 15'h6591: d <= 8'h33; 15'h6592: d <= 8'h37; 15'h6593: d <= 8'h3B;
                15'h6594: d <= 8'h44; 15'h6595: d <= 8'h48; 15'h6596: d <= 8'h4C; 15'h6597: d <= 8'h41;
                15'h6598: d <= 8'h49; 15'h6599: d <= 8'h4D; 15'h659A: d <= 8'h42; 15'h659B: d <= 8'h46;
                15'h659C: d <= 8'h4E; 15'h659D: d <= 8'h43; 15'h659E: d <= 8'h47; 15'h659F: d <= 8'h4B;
                15'h65A0: d <= 8'h50; 15'h65A1: d <= 8'h55; 15'h65A2: d <= 8'h5A; 15'h65A3: d <= 8'h5F;
                15'h65A4: d <= 8'h60; 15'h65A5: d <= 8'h65; 15'h65A6: d <= 8'h6A; 15'h65A7: d <= 8'h6F;
                15'h65A8: d <= 8'h74; 15'h65A9: d <= 8'h78; 15'h65AA: d <= 8'h7C; 15'h65AB: d <= 8'h71;
                15'h65AC: d <= 8'h79; 15'h65AD: d <= 8'h7D; 15'h65AE: d <= 8'h72; 15'h65AF: d <= 8'h76;
                15'h65B0: d <= 8'h7E; 15'h65B1: d <= 8'h73; 15'h65B2: d <= 8'h77; 15'h65B3: d <= 8'h7B;
                15'h65B4: d <= 8'h84; 15'h65B5: d <= 8'h88; 15'h65B6: d <= 8'h8C; 15'h65B7: d <= 8'h81;
                15'h65B8: d <= 8'h89; 15'h65B9: d <= 8'h8D; 15'h65BA: d <= 8'h82; 15'h65BB: d <= 8'h86;
                15'h65BC: d <= 8'h8E; 15'h65BD: d <= 8'h83; 15'h65BE: d <= 8'h87; 15'h65BF: d <= 8'h8B;
                15'h65C0: d <= 8'h90; 15'h65C1: d <= 8'h95; 15'h65C2: d <= 8'h9A; 15'h65C3: d <= 8'h9F;
                15'h65C4: d <= 8'hA4; 15'h65C5: d <= 8'hA8; 15'h65C6: d <= 8'hAC; 15'h65C7: d <= 8'hA1;
                15'h65C8: d <= 8'hA9; 15'h65C9: d <= 8'hAD; 15'h65CA: d <= 8'hA2; 15'h65CB: d <= 8'hA6;
                15'h65CC: d <= 8'hAE; 15'h65CD: d <= 8'hA3; 15'h65CE: d <= 8'hA7; 15'h65CF: d <= 8'hAB;
                15'h65D0: d <= 8'hB4; 15'h65D1: d <= 8'hB8; 15'h65D2: d <= 8'hBC; 15'h65D3: d <= 8'hB1;
                15'h65D4: d <= 8'hB9; 15'h65D5: d <= 8'hBD; 15'h65D6: d <= 8'hB2; 15'h65D7: d <= 8'hB6;
                15'h65D8: d <= 8'hBE; 15'h65D9: d <= 8'hB3; 15'h65DA: d <= 8'hB7; 15'h65DB: d <= 8'hBB;
                15'h65DC: d <= 8'hC4; 15'h65DD: d <= 8'hC8; 15'h65DE: d <= 8'hCC; 15'h65DF: d <= 8'hC1;
                15'h65E0: d <= 8'hC9; 15'h65E1: d <= 8'hCD; 15'h65E2: d <= 8'hC2; 15'h65E3: d <= 8'hC6;
                15'h65E4: d <= 8'hCE; 15'h65E5: d <= 8'hC3; 15'h65E6: d <= 8'hC7; 15'h65E7: d <= 8'hCB;
                15'h65E8: d <= 8'hC0; 15'h65E9: d <= 8'hC5; 15'h65EA: d <= 8'hCA; 15'h65EB: d <= 8'hCF;
                15'h65EC: d <= 8'hD0; 15'h65ED: d <= 8'hD5; 15'h65EE: d <= 8'hDA; 15'h65EF: d <= 8'hDF;
                15'h65F0: d <= 8'h74; 15'h65F1: d <= 8'h78; 15'h65F2: d <= 8'h7C; 15'h65F3: d <= 8'h71;
                15'h65F4: d <= 8'h79; 15'h65F5: d <= 8'h7D; 15'h65F6: d <= 8'h72; 15'h65F7: d <= 8'h76;
                15'h65F8: d <= 8'h7E; 15'h65F9: d <= 8'h73; 15'h65FA: d <= 8'h77; 15'h65FB: d <= 8'h7B;
                15'h65FC: d <= 8'hA0; 15'h65FD: d <= 8'hA5; 15'h65FE: d <= 8'hAA; 15'h65FF: d <= 8'hAF;
                15'h6600: d <= 8'h00; 15'h6601: d <= 8'h00; 15'h6602: d <= 8'h00; 15'h6603: d <= 8'h00;
                15'h6604: d <= 8'h00; 15'h6605: d <= 8'h00; 15'h6606: d <= 8'h00; 15'h6607: d <= 8'h00;
                15'h6608: d <= 8'h00; 15'h6609: d <= 8'h00; 15'h660A: d <= 8'h00; 15'h660B: d <= 8'h00;
                15'h660C: d <= 8'h00; 15'h660D: d <= 8'h00; 15'h660E: d <= 8'h00; 15'h660F: d <= 8'h00;
                15'h6610: d <= 8'h00; 15'h6611: d <= 8'h00; 15'h6612: d <= 8'h00; 15'h6613: d <= 8'h00;
                15'h6614: d <= 8'h00; 15'h6615: d <= 8'h00; 15'h6616: d <= 8'h00; 15'h6617: d <= 8'h00;
                15'h6618: d <= 8'h00; 15'h6619: d <= 8'h00; 15'h661A: d <= 8'h00; 15'h661B: d <= 8'h00;
                15'h661C: d <= 8'h00; 15'h661D: d <= 8'h00; 15'h661E: d <= 8'h00; 15'h661F: d <= 8'h00;
                15'h6620: d <= 8'h00; 15'h6621: d <= 8'h00; 15'h6622: d <= 8'h00; 15'h6623: d <= 8'h00;
                15'h6624: d <= 8'h00; 15'h6625: d <= 8'h00; 15'h6626: d <= 8'h00; 15'h6627: d <= 8'h00;
                15'h6628: d <= 8'h00; 15'h6629: d <= 8'h00; 15'h662A: d <= 8'h00; 15'h662B: d <= 8'h00;
                15'h662C: d <= 8'h00; 15'h662D: d <= 8'h00; 15'h662E: d <= 8'h00; 15'h662F: d <= 8'hAF;
                15'h6630: d <= 8'h00; 15'h6631: d <= 8'h00; 15'h6632: d <= 8'h00; 15'h6633: d <= 8'h00;
                15'h6634: d <= 8'h00; 15'h6635: d <= 8'h00; 15'h6636: d <= 8'h00; 15'h6637: d <= 8'h00;
                15'h6638: d <= 8'h00; 15'h6639: d <= 8'h00; 15'h663A: d <= 8'h00; 15'h663B: d <= 8'h00;
                15'h663C: d <= 8'h00; 15'h663D: d <= 8'h00; 15'h663E: d <= 8'h00; 15'h663F: d <= 8'h00;
                15'h6640: d <= 8'h00; 15'h6641: d <= 8'h00; 15'h6642: d <= 8'h00; 15'h6643: d <= 8'h00;
                15'h6644: d <= 8'h00; 15'h6645: d <= 8'h00; 15'h6646: d <= 8'h00; 15'h6647: d <= 8'h00;
                15'h6648: d <= 8'h00; 15'h6649: d <= 8'h00; 15'h664A: d <= 8'h00; 15'h664B: d <= 8'h00;
                15'h664C: d <= 8'h00; 15'h664D: d <= 8'h00; 15'h664E: d <= 8'h00; 15'h664F: d <= 8'h00;
                15'h6650: d <= 8'h00; 15'h6651: d <= 8'h00; 15'h6652: d <= 8'h00; 15'h6653: d <= 8'h00;
                15'h6654: d <= 8'h00; 15'h6655: d <= 8'h00; 15'h6656: d <= 8'h00; 15'h6657: d <= 8'h00;
                15'h6658: d <= 8'h45; 15'h6659: d <= 8'h35; 15'h665A: d <= 8'hAA; 15'h665B: d <= 8'h00;
                15'h665C: d <= 8'h00; 15'h665D: d <= 8'h00; 15'h665E: d <= 8'h00; 15'h665F: d <= 8'h00;
                15'h6660: d <= 8'h00; 15'h6661: d <= 8'h00; 15'h6662: d <= 8'h00; 15'h6663: d <= 8'h00;
                15'h6664: d <= 8'h00; 15'h6665: d <= 8'h00; 15'h6666: d <= 8'h00; 15'h6667: d <= 8'h00;
                15'h6668: d <= 8'h00; 15'h6669: d <= 8'h00; 15'h666A: d <= 8'h00; 15'h666B: d <= 8'h00;
                15'h666C: d <= 8'h00; 15'h666D: d <= 8'h00; 15'h666E: d <= 8'h00; 15'h666F: d <= 8'h00;
                15'h6670: d <= 8'h00; 15'h6671: d <= 8'h00; 15'h6672: d <= 8'h00; 15'h6673: d <= 8'h00;
                15'h6674: d <= 8'h00; 15'h6675: d <= 8'h00; 15'h6676: d <= 8'h00; 15'h6677: d <= 8'h00;
                15'h6678: d <= 8'h00; 15'h6679: d <= 8'h00; 15'h667A: d <= 8'h00; 15'h667B: d <= 8'h00;
                15'h667C: d <= 8'h00; 15'h667D: d <= 8'h00; 15'h667E: d <= 8'h00; 15'h667F: d <= 8'hE0;
                15'h6680: d <= 8'h10; 15'h6681: d <= 8'h15; 15'h6682: d <= 8'h1A; 15'h6683: d <= 8'h1F;
                15'h6684: d <= 8'h20; 15'h6685: d <= 8'h25; 15'h6686: d <= 8'h2A; 15'h6687: d <= 8'h2F;
                15'h6688: d <= 8'h34; 15'h6689: d <= 8'h38; 15'h668A: d <= 8'h3C; 15'h668B: d <= 8'h31;
                15'h668C: d <= 8'h39; 15'h668D: d <= 8'h3D; 15'h668E: d <= 8'h32; 15'h668F: d <= 8'h36;
                15'h6690: d <= 8'h3E; 15'h6691: d <= 8'h33; 15'h6692: d <= 8'h37; 15'h6693: d <= 8'h3B;
                15'h6694: d <= 8'h44; 15'h6695: d <= 8'h48; 15'h6696: d <= 8'h4C; 15'h6697: d <= 8'h41;
                15'h6698: d <= 8'h49; 15'h6699: d <= 8'h4D; 15'h669A: d <= 8'h42; 15'h669B: d <= 8'h46;
                15'h669C: d <= 8'h4E; 15'h669D: d <= 8'h43; 15'h669E: d <= 8'h47; 15'h669F: d <= 8'h4B;
                15'h66A0: d <= 8'h50; 15'h66A1: d <= 8'h55; 15'h66A2: d <= 8'h5A; 15'h66A3: d <= 8'h5F;
                15'h66A4: d <= 8'h60; 15'h66A5: d <= 8'h65; 15'h66A6: d <= 8'h6A; 15'h66A7: d <= 8'h6F;
                15'h66A8: d <= 8'h74; 15'h66A9: d <= 8'h78; 15'h66AA: d <= 8'h7C; 15'h66AB: d <= 8'h71;
                15'h66AC: d <= 8'h79; 15'h66AD: d <= 8'h7D; 15'h66AE: d <= 8'h72; 15'h66AF: d <= 8'h76;
                15'h66B0: d <= 8'h7E; 15'h66B1: d <= 8'h73; 15'h66B2: d <= 8'h77; 15'h66B3: d <= 8'h7B;
                15'h66B4: d <= 8'h84; 15'h66B5: d <= 8'h88; 15'h66B6: d <= 8'h8C; 15'h66B7: d <= 8'h81;
                15'h66B8: d <= 8'h89; 15'h66B9: d <= 8'h8D; 15'h66BA: d <= 8'h82; 15'h66BB: d <= 8'h86;
                15'h66BC: d <= 8'h8E; 15'h66BD: d <= 8'h83; 15'h66BE: d <= 8'h87; 15'h66BF: d <= 8'h8B;
                15'h66C0: d <= 8'h90; 15'h66C1: d <= 8'h95; 15'h66C2: d <= 8'h9A; 15'h66C3: d <= 8'h9F;
                15'h66C4: d <= 8'hA4; 15'h66C5: d <= 8'hA8; 15'h66C6: d <= 8'hAC; 15'h66C7: d <= 8'hA1;
                15'h66C8: d <= 8'hA9; 15'h66C9: d <= 8'hAD; 15'h66CA: d <= 8'hA2; 15'h66CB: d <= 8'hA6;
                15'h66CC: d <= 8'hAE; 15'h66CD: d <= 8'hA3; 15'h66CE: d <= 8'hA7; 15'h66CF: d <= 8'hAB;
                15'h66D0: d <= 8'hB4; 15'h66D1: d <= 8'hB8; 15'h66D2: d <= 8'hBC; 15'h66D3: d <= 8'hB1;
                15'h66D4: d <= 8'hB9; 15'h66D5: d <= 8'hBD; 15'h66D6: d <= 8'hB2; 15'h66D7: d <= 8'hB6;
                15'h66D8: d <= 8'hBE; 15'h66D9: d <= 8'hB3; 15'h66DA: d <= 8'hB7; 15'h66DB: d <= 8'hBB;
                15'h66DC: d <= 8'hC4; 15'h66DD: d <= 8'hC8; 15'h66DE: d <= 8'hCC; 15'h66DF: d <= 8'hC1;
                15'h66E0: d <= 8'hC9; 15'h66E1: d <= 8'hCD; 15'h66E2: d <= 8'hC2; 15'h66E3: d <= 8'hC6;
                15'h66E4: d <= 8'hCE; 15'h66E5: d <= 8'hC3; 15'h66E6: d <= 8'hC7; 15'h66E7: d <= 8'hCB;
                15'h66E8: d <= 8'hC0; 15'h66E9: d <= 8'hC5; 15'h66EA: d <= 8'hCA; 15'h66EB: d <= 8'hCF;
                15'h66EC: d <= 8'hD0; 15'h66ED: d <= 8'hD5; 15'h66EE: d <= 8'hDA; 15'h66EF: d <= 8'hDF;
                15'h66F0: d <= 8'h74; 15'h66F1: d <= 8'h78; 15'h66F2: d <= 8'h7C; 15'h66F3: d <= 8'h71;
                15'h66F4: d <= 8'h79; 15'h66F5: d <= 8'h7D; 15'h66F6: d <= 8'h72; 15'h66F7: d <= 8'h76;
                15'h66F8: d <= 8'h7E; 15'h66F9: d <= 8'h73; 15'h66FA: d <= 8'h77; 15'h66FB: d <= 8'h7B;
                15'h66FC: d <= 8'hA0; 15'h66FD: d <= 8'hA5; 15'h66FE: d <= 8'hAA; 15'h66FF: d <= 8'hAF;
                15'h6700: d <= 8'h00; 15'h6701: d <= 8'h00; 15'h6702: d <= 8'h00; 15'h6703: d <= 8'h00;
                15'h6704: d <= 8'h00; 15'h6705: d <= 8'h00; 15'h6706: d <= 8'h00; 15'h6707: d <= 8'h00;
                15'h6708: d <= 8'h00; 15'h6709: d <= 8'h00; 15'h670A: d <= 8'h00; 15'h670B: d <= 8'h00;
                15'h670C: d <= 8'h00; 15'h670D: d <= 8'h00; 15'h670E: d <= 8'h00; 15'h670F: d <= 8'h00;
                15'h6710: d <= 8'h00; 15'h6711: d <= 8'h00; 15'h6712: d <= 8'h00; 15'h6713: d <= 8'h00;
                15'h6714: d <= 8'h00; 15'h6715: d <= 8'h00; 15'h6716: d <= 8'h00; 15'h6717: d <= 8'h00;
                15'h6718: d <= 8'h00; 15'h6719: d <= 8'h00; 15'h671A: d <= 8'h00; 15'h671B: d <= 8'h00;
                15'h671C: d <= 8'h00; 15'h671D: d <= 8'h00; 15'h671E: d <= 8'h00; 15'h671F: d <= 8'h00;
                15'h6720: d <= 8'h00; 15'h6721: d <= 8'h00; 15'h6722: d <= 8'h00; 15'h6723: d <= 8'h00;
                15'h6724: d <= 8'h00; 15'h6725: d <= 8'h00; 15'h6726: d <= 8'h00; 15'h6727: d <= 8'h00;
                15'h6728: d <= 8'h00; 15'h6729: d <= 8'h00; 15'h672A: d <= 8'h00; 15'h672B: d <= 8'h00;
                15'h672C: d <= 8'h00; 15'h672D: d <= 8'h00; 15'h672E: d <= 8'h00; 15'h672F: d <= 8'hAF;
                15'h6730: d <= 8'h00; 15'h6731: d <= 8'h00; 15'h6732: d <= 8'h00; 15'h6733: d <= 8'h00;
                15'h6734: d <= 8'h00; 15'h6735: d <= 8'h00; 15'h6736: d <= 8'h00; 15'h6737: d <= 8'h00;
                15'h6738: d <= 8'h00; 15'h6739: d <= 8'h00; 15'h673A: d <= 8'h00; 15'h673B: d <= 8'h00;
                15'h673C: d <= 8'h00; 15'h673D: d <= 8'h00; 15'h673E: d <= 8'h00; 15'h673F: d <= 8'h00;
                15'h6740: d <= 8'h00; 15'h6741: d <= 8'h00; 15'h6742: d <= 8'h00; 15'h6743: d <= 8'h00;
                15'h6744: d <= 8'h00; 15'h6745: d <= 8'h00; 15'h6746: d <= 8'h00; 15'h6747: d <= 8'h00;
                15'h6748: d <= 8'h00; 15'h6749: d <= 8'h00; 15'h674A: d <= 8'h00; 15'h674B: d <= 8'h00;
                15'h674C: d <= 8'h00; 15'h674D: d <= 8'h00; 15'h674E: d <= 8'h00; 15'h674F: d <= 8'h00;
                15'h6750: d <= 8'h00; 15'h6751: d <= 8'h00; 15'h6752: d <= 8'h00; 15'h6753: d <= 8'h00;
                15'h6754: d <= 8'h00; 15'h6755: d <= 8'h00; 15'h6756: d <= 8'h00; 15'h6757: d <= 8'h00;
                15'h6758: d <= 8'h45; 15'h6759: d <= 8'h35; 15'h675A: d <= 8'hAA; 15'h675B: d <= 8'h00;
                15'h675C: d <= 8'h00; 15'h675D: d <= 8'h00; 15'h675E: d <= 8'h00; 15'h675F: d <= 8'h00;
                15'h6760: d <= 8'h00; 15'h6761: d <= 8'h00; 15'h6762: d <= 8'h00; 15'h6763: d <= 8'h00;
                15'h6764: d <= 8'h00; 15'h6765: d <= 8'h00; 15'h6766: d <= 8'h00; 15'h6767: d <= 8'h00;
                15'h6768: d <= 8'h00; 15'h6769: d <= 8'h00; 15'h676A: d <= 8'h00; 15'h676B: d <= 8'h00;
                15'h676C: d <= 8'h00; 15'h676D: d <= 8'h00; 15'h676E: d <= 8'h00; 15'h676F: d <= 8'h00;
                15'h6770: d <= 8'h00; 15'h6771: d <= 8'h00; 15'h6772: d <= 8'h00; 15'h6773: d <= 8'h00;
                15'h6774: d <= 8'h00; 15'h6775: d <= 8'h00; 15'h6776: d <= 8'h00; 15'h6777: d <= 8'h00;
                15'h6778: d <= 8'h00; 15'h6779: d <= 8'h00; 15'h677A: d <= 8'h00; 15'h677B: d <= 8'h00;
                15'h677C: d <= 8'h00; 15'h677D: d <= 8'h00; 15'h677E: d <= 8'h00; 15'h677F: d <= 8'hE0;
                15'h6780: d <= 8'h10; 15'h6781: d <= 8'h15; 15'h6782: d <= 8'h1A; 15'h6783: d <= 8'h1F;
                15'h6784: d <= 8'h20; 15'h6785: d <= 8'h25; 15'h6786: d <= 8'h2A; 15'h6787: d <= 8'h2F;
                15'h6788: d <= 8'h34; 15'h6789: d <= 8'h38; 15'h678A: d <= 8'h3C; 15'h678B: d <= 8'h31;
                15'h678C: d <= 8'h39; 15'h678D: d <= 8'h3D; 15'h678E: d <= 8'h32; 15'h678F: d <= 8'h36;
                15'h6790: d <= 8'h3E; 15'h6791: d <= 8'h33; 15'h6792: d <= 8'h37; 15'h6793: d <= 8'h3B;
                15'h6794: d <= 8'h44; 15'h6795: d <= 8'h48; 15'h6796: d <= 8'h4C; 15'h6797: d <= 8'h41;
                15'h6798: d <= 8'h49; 15'h6799: d <= 8'h4D; 15'h679A: d <= 8'h42; 15'h679B: d <= 8'h46;
                15'h679C: d <= 8'h4E; 15'h679D: d <= 8'h43; 15'h679E: d <= 8'h47; 15'h679F: d <= 8'h4B;
                15'h67A0: d <= 8'h50; 15'h67A1: d <= 8'h55; 15'h67A2: d <= 8'h5A; 15'h67A3: d <= 8'h5F;
                15'h67A4: d <= 8'h60; 15'h67A5: d <= 8'h65; 15'h67A6: d <= 8'h6A; 15'h67A7: d <= 8'h6F;
                15'h67A8: d <= 8'h74; 15'h67A9: d <= 8'h78; 15'h67AA: d <= 8'h7C; 15'h67AB: d <= 8'h71;
                15'h67AC: d <= 8'h79; 15'h67AD: d <= 8'h7D; 15'h67AE: d <= 8'h72; 15'h67AF: d <= 8'h76;
                15'h67B0: d <= 8'h7E; 15'h67B1: d <= 8'h73; 15'h67B2: d <= 8'h77; 15'h67B3: d <= 8'h7B;
                15'h67B4: d <= 8'h84; 15'h67B5: d <= 8'h88; 15'h67B6: d <= 8'h8C; 15'h67B7: d <= 8'h81;
                15'h67B8: d <= 8'h89; 15'h67B9: d <= 8'h8D; 15'h67BA: d <= 8'h82; 15'h67BB: d <= 8'h86;
                15'h67BC: d <= 8'h8E; 15'h67BD: d <= 8'h83; 15'h67BE: d <= 8'h87; 15'h67BF: d <= 8'h8B;
                15'h67C0: d <= 8'h90; 15'h67C1: d <= 8'h95; 15'h67C2: d <= 8'h9A; 15'h67C3: d <= 8'h9F;
                15'h67C4: d <= 8'hA4; 15'h67C5: d <= 8'hA8; 15'h67C6: d <= 8'hAC; 15'h67C7: d <= 8'hA1;
                15'h67C8: d <= 8'hA9; 15'h67C9: d <= 8'hAD; 15'h67CA: d <= 8'hA2; 15'h67CB: d <= 8'hA6;
                15'h67CC: d <= 8'hAE; 15'h67CD: d <= 8'hA3; 15'h67CE: d <= 8'hA7; 15'h67CF: d <= 8'hAB;
                15'h67D0: d <= 8'hB4; 15'h67D1: d <= 8'hB8; 15'h67D2: d <= 8'hBC; 15'h67D3: d <= 8'hB1;
                15'h67D4: d <= 8'hB9; 15'h67D5: d <= 8'hBD; 15'h67D6: d <= 8'hB2; 15'h67D7: d <= 8'hB6;
                15'h67D8: d <= 8'hBE; 15'h67D9: d <= 8'hB3; 15'h67DA: d <= 8'hB7; 15'h67DB: d <= 8'hBB;
                15'h67DC: d <= 8'hC4; 15'h67DD: d <= 8'hC8; 15'h67DE: d <= 8'hCC; 15'h67DF: d <= 8'hC1;
                15'h67E0: d <= 8'hC9; 15'h67E1: d <= 8'hCD; 15'h67E2: d <= 8'hC2; 15'h67E3: d <= 8'hC6;
                15'h67E4: d <= 8'hCE; 15'h67E5: d <= 8'hC3; 15'h67E6: d <= 8'hC7; 15'h67E7: d <= 8'hCB;
                15'h67E8: d <= 8'hC0; 15'h67E9: d <= 8'hC5; 15'h67EA: d <= 8'hCA; 15'h67EB: d <= 8'hCF;
                15'h67EC: d <= 8'hD0; 15'h67ED: d <= 8'hD5; 15'h67EE: d <= 8'hDA; 15'h67EF: d <= 8'hDF;
                15'h67F0: d <= 8'h74; 15'h67F1: d <= 8'h78; 15'h67F2: d <= 8'h7C; 15'h67F3: d <= 8'h71;
                15'h67F4: d <= 8'h79; 15'h67F5: d <= 8'h7D; 15'h67F6: d <= 8'h72; 15'h67F7: d <= 8'h76;
                15'h67F8: d <= 8'h7E; 15'h67F9: d <= 8'h73; 15'h67FA: d <= 8'h77; 15'h67FB: d <= 8'h7B;
                15'h67FC: d <= 8'hA0; 15'h67FD: d <= 8'hA5; 15'h67FE: d <= 8'hAA; 15'h67FF: d <= 8'hAF;
                15'h6800: d <= 8'h00; 15'h6801: d <= 8'h00; 15'h6802: d <= 8'h00; 15'h6803: d <= 8'h00;
                15'h6804: d <= 8'h00; 15'h6805: d <= 8'h00; 15'h6806: d <= 8'h00; 15'h6807: d <= 8'h00;
                15'h6808: d <= 8'h00; 15'h6809: d <= 8'h00; 15'h680A: d <= 8'h00; 15'h680B: d <= 8'h00;
                15'h680C: d <= 8'h00; 15'h680D: d <= 8'h00; 15'h680E: d <= 8'h00; 15'h680F: d <= 8'h00;
                15'h6810: d <= 8'h00; 15'h6811: d <= 8'h00; 15'h6812: d <= 8'h00; 15'h6813: d <= 8'h00;
                15'h6814: d <= 8'h00; 15'h6815: d <= 8'h00; 15'h6816: d <= 8'h00; 15'h6817: d <= 8'h00;
                15'h6818: d <= 8'h00; 15'h6819: d <= 8'h00; 15'h681A: d <= 8'h00; 15'h681B: d <= 8'h00;
                15'h681C: d <= 8'h00; 15'h681D: d <= 8'h00; 15'h681E: d <= 8'h00; 15'h681F: d <= 8'h00;
                15'h6820: d <= 8'h00; 15'h6821: d <= 8'h00; 15'h6822: d <= 8'h00; 15'h6823: d <= 8'h00;
                15'h6824: d <= 8'h00; 15'h6825: d <= 8'h00; 15'h6826: d <= 8'h00; 15'h6827: d <= 8'h00;
                15'h6828: d <= 8'h00; 15'h6829: d <= 8'h00; 15'h682A: d <= 8'h00; 15'h682B: d <= 8'h00;
                15'h682C: d <= 8'h00; 15'h682D: d <= 8'h00; 15'h682E: d <= 8'h00; 15'h682F: d <= 8'h7B;
                15'h6830: d <= 8'h00; 15'h6831: d <= 8'h00; 15'h6832: d <= 8'h00; 15'h6833: d <= 8'h00;
                15'h6834: d <= 8'h00; 15'h6835: d <= 8'h00; 15'h6836: d <= 8'h00; 15'h6837: d <= 8'h00;
                15'h6838: d <= 8'h00; 15'h6839: d <= 8'h00; 15'h683A: d <= 8'h00; 15'h683B: d <= 8'h00;
                15'h683C: d <= 8'h00; 15'h683D: d <= 8'h00; 15'h683E: d <= 8'h00; 15'h683F: d <= 8'h00;
                15'h6840: d <= 8'h00; 15'h6841: d <= 8'h00; 15'h6842: d <= 8'h00; 15'h6843: d <= 8'h00;
                15'h6844: d <= 8'h00; 15'h6845: d <= 8'h00; 15'h6846: d <= 8'h00; 15'h6847: d <= 8'h00;
                15'h6848: d <= 8'h00; 15'h6849: d <= 8'h00; 15'h684A: d <= 8'h00; 15'h684B: d <= 8'h00;
                15'h684C: d <= 8'h00; 15'h684D: d <= 8'h00; 15'h684E: d <= 8'h00; 15'h684F: d <= 8'h00;
                15'h6850: d <= 8'h00; 15'h6851: d <= 8'h00; 15'h6852: d <= 8'h00; 15'h6853: d <= 8'h00;
                15'h6854: d <= 8'h00; 15'h6855: d <= 8'h00; 15'h6856: d <= 8'h00; 15'h6857: d <= 8'h00;
                15'h6858: d <= 8'h45; 15'h6859: d <= 8'h35; 15'h685A: d <= 8'h32; 15'h685B: d <= 8'h00;
                15'h685C: d <= 8'h00; 15'h685D: d <= 8'h00; 15'h685E: d <= 8'h00; 15'h685F: d <= 8'h00;
                15'h6860: d <= 8'h00; 15'h6861: d <= 8'h00; 15'h6862: d <= 8'h00; 15'h6863: d <= 8'h00;
                15'h6864: d <= 8'h00; 15'h6865: d <= 8'h00; 15'h6866: d <= 8'h00; 15'h6867: d <= 8'h00;
                15'h6868: d <= 8'h00; 15'h6869: d <= 8'h00; 15'h686A: d <= 8'h00; 15'h686B: d <= 8'h00;
                15'h686C: d <= 8'h00; 15'h686D: d <= 8'h00; 15'h686E: d <= 8'h00; 15'h686F: d <= 8'h00;
                15'h6870: d <= 8'h00; 15'h6871: d <= 8'h00; 15'h6872: d <= 8'h00; 15'h6873: d <= 8'h00;
                15'h6874: d <= 8'h00; 15'h6875: d <= 8'h00; 15'h6876: d <= 8'h00; 15'h6877: d <= 8'h00;
                15'h6878: d <= 8'h00; 15'h6879: d <= 8'h00; 15'h687A: d <= 8'h00; 15'h687B: d <= 8'h00;
                15'h687C: d <= 8'h00; 15'h687D: d <= 8'h00; 15'h687E: d <= 8'h00; 15'h687F: d <= 8'hE0;
                15'h6880: d <= 8'h10; 15'h6881: d <= 8'h15; 15'h6882: d <= 8'h1A; 15'h6883: d <= 8'h1F;
                15'h6884: d <= 8'h20; 15'h6885: d <= 8'h25; 15'h6886: d <= 8'h2A; 15'h6887: d <= 8'h2F;
                15'h6888: d <= 8'h34; 15'h6889: d <= 8'h38; 15'h688A: d <= 8'h3C; 15'h688B: d <= 8'h31;
                15'h688C: d <= 8'h39; 15'h688D: d <= 8'h3D; 15'h688E: d <= 8'h32; 15'h688F: d <= 8'h36;
                15'h6890: d <= 8'h3E; 15'h6891: d <= 8'h33; 15'h6892: d <= 8'h37; 15'h6893: d <= 8'h3B;
                15'h6894: d <= 8'h44; 15'h6895: d <= 8'h48; 15'h6896: d <= 8'h4C; 15'h6897: d <= 8'h41;
                15'h6898: d <= 8'h49; 15'h6899: d <= 8'h4D; 15'h689A: d <= 8'h42; 15'h689B: d <= 8'h46;
                15'h689C: d <= 8'h4E; 15'h689D: d <= 8'h43; 15'h689E: d <= 8'h47; 15'h689F: d <= 8'h4B;
                15'h68A0: d <= 8'h50; 15'h68A1: d <= 8'h55; 15'h68A2: d <= 8'h5A; 15'h68A3: d <= 8'h5F;
                15'h68A4: d <= 8'h60; 15'h68A5: d <= 8'h65; 15'h68A6: d <= 8'h6A; 15'h68A7: d <= 8'h6F;
                15'h68A8: d <= 8'h74; 15'h68A9: d <= 8'h78; 15'h68AA: d <= 8'h7C; 15'h68AB: d <= 8'h71;
                15'h68AC: d <= 8'h79; 15'h68AD: d <= 8'h7D; 15'h68AE: d <= 8'h72; 15'h68AF: d <= 8'h76;
                15'h68B0: d <= 8'h7E; 15'h68B1: d <= 8'h73; 15'h68B2: d <= 8'h77; 15'h68B3: d <= 8'h7B;
                15'h68B4: d <= 8'h84; 15'h68B5: d <= 8'h88; 15'h68B6: d <= 8'h8C; 15'h68B7: d <= 8'h81;
                15'h68B8: d <= 8'h89; 15'h68B9: d <= 8'h8D; 15'h68BA: d <= 8'h82; 15'h68BB: d <= 8'h86;
                15'h68BC: d <= 8'h8E; 15'h68BD: d <= 8'h83; 15'h68BE: d <= 8'h87; 15'h68BF: d <= 8'h8B;
                15'h68C0: d <= 8'h90; 15'h68C1: d <= 8'h95; 15'h68C2: d <= 8'h9A; 15'h68C3: d <= 8'h9F;
                15'h68C4: d <= 8'hA4; 15'h68C5: d <= 8'hA8; 15'h68C6: d <= 8'hAC; 15'h68C7: d <= 8'hA1;
                15'h68C8: d <= 8'hA9; 15'h68C9: d <= 8'hAD; 15'h68CA: d <= 8'hA2; 15'h68CB: d <= 8'hA6;
                15'h68CC: d <= 8'hAE; 15'h68CD: d <= 8'hA3; 15'h68CE: d <= 8'hA7; 15'h68CF: d <= 8'hAB;
                15'h68D0: d <= 8'hB4; 15'h68D1: d <= 8'hB8; 15'h68D2: d <= 8'hBC; 15'h68D3: d <= 8'hB1;
                15'h68D4: d <= 8'hB9; 15'h68D5: d <= 8'hBD; 15'h68D6: d <= 8'hB2; 15'h68D7: d <= 8'hB6;
                15'h68D8: d <= 8'hBE; 15'h68D9: d <= 8'hB3; 15'h68DA: d <= 8'hB7; 15'h68DB: d <= 8'hBB;
                15'h68DC: d <= 8'hC4; 15'h68DD: d <= 8'hC8; 15'h68DE: d <= 8'hCC; 15'h68DF: d <= 8'hC1;
                15'h68E0: d <= 8'hC9; 15'h68E1: d <= 8'hCD; 15'h68E2: d <= 8'hC2; 15'h68E3: d <= 8'hC6;
                15'h68E4: d <= 8'hCE; 15'h68E5: d <= 8'hC3; 15'h68E6: d <= 8'hC7; 15'h68E7: d <= 8'hCB;
                15'h68E8: d <= 8'hC0; 15'h68E9: d <= 8'hC5; 15'h68EA: d <= 8'hCA; 15'h68EB: d <= 8'hCF;
                15'h68EC: d <= 8'hD0; 15'h68ED: d <= 8'hD5; 15'h68EE: d <= 8'hDA; 15'h68EF: d <= 8'hDF;
                15'h68F0: d <= 8'h74; 15'h68F1: d <= 8'h78; 15'h68F2: d <= 8'h7C; 15'h68F3: d <= 8'h71;
                15'h68F4: d <= 8'h79; 15'h68F5: d <= 8'h7D; 15'h68F6: d <= 8'h72; 15'h68F7: d <= 8'h76;
                15'h68F8: d <= 8'h7E; 15'h68F9: d <= 8'h73; 15'h68FA: d <= 8'h77; 15'h68FB: d <= 8'h7B;
                15'h68FC: d <= 8'hA0; 15'h68FD: d <= 8'hA5; 15'h68FE: d <= 8'hAA; 15'h68FF: d <= 8'hAF;
                15'h6900: d <= 8'h00; 15'h6901: d <= 8'h00; 15'h6902: d <= 8'h00; 15'h6903: d <= 8'h00;
                15'h6904: d <= 8'h00; 15'h6905: d <= 8'h00; 15'h6906: d <= 8'h00; 15'h6907: d <= 8'h00;
                15'h6908: d <= 8'h00; 15'h6909: d <= 8'h00; 15'h690A: d <= 8'h00; 15'h690B: d <= 8'h00;
                15'h690C: d <= 8'h00; 15'h690D: d <= 8'h00; 15'h690E: d <= 8'h00; 15'h690F: d <= 8'h00;
                15'h6910: d <= 8'h00; 15'h6911: d <= 8'h00; 15'h6912: d <= 8'h00; 15'h6913: d <= 8'h00;
                15'h6914: d <= 8'h00; 15'h6915: d <= 8'h00; 15'h6916: d <= 8'h00; 15'h6917: d <= 8'h00;
                15'h6918: d <= 8'h00; 15'h6919: d <= 8'h00; 15'h691A: d <= 8'h00; 15'h691B: d <= 8'h00;
                15'h691C: d <= 8'h00; 15'h691D: d <= 8'h00; 15'h691E: d <= 8'h00; 15'h691F: d <= 8'h00;
                15'h6920: d <= 8'h00; 15'h6921: d <= 8'h00; 15'h6922: d <= 8'h00; 15'h6923: d <= 8'h00;
                15'h6924: d <= 8'h00; 15'h6925: d <= 8'h00; 15'h6926: d <= 8'h00; 15'h6927: d <= 8'h00;
                15'h6928: d <= 8'h00; 15'h6929: d <= 8'h00; 15'h692A: d <= 8'h00; 15'h692B: d <= 8'h00;
                15'h692C: d <= 8'h00; 15'h692D: d <= 8'h00; 15'h692E: d <= 8'h00; 15'h692F: d <= 8'h7B;
                15'h6930: d <= 8'h00; 15'h6931: d <= 8'h00; 15'h6932: d <= 8'h00; 15'h6933: d <= 8'h00;
                15'h6934: d <= 8'h00; 15'h6935: d <= 8'h00; 15'h6936: d <= 8'h00; 15'h6937: d <= 8'h00;
                15'h6938: d <= 8'h00; 15'h6939: d <= 8'h00; 15'h693A: d <= 8'h00; 15'h693B: d <= 8'h00;
                15'h693C: d <= 8'h00; 15'h693D: d <= 8'h00; 15'h693E: d <= 8'h00; 15'h693F: d <= 8'h00;
                15'h6940: d <= 8'h00; 15'h6941: d <= 8'h00; 15'h6942: d <= 8'h00; 15'h6943: d <= 8'h00;
                15'h6944: d <= 8'h00; 15'h6945: d <= 8'h00; 15'h6946: d <= 8'h00; 15'h6947: d <= 8'h00;
                15'h6948: d <= 8'h00; 15'h6949: d <= 8'h00; 15'h694A: d <= 8'h00; 15'h694B: d <= 8'h00;
                15'h694C: d <= 8'h00; 15'h694D: d <= 8'h00; 15'h694E: d <= 8'h00; 15'h694F: d <= 8'h00;
                15'h6950: d <= 8'h00; 15'h6951: d <= 8'h00; 15'h6952: d <= 8'h00; 15'h6953: d <= 8'h00;
                15'h6954: d <= 8'h00; 15'h6955: d <= 8'h00; 15'h6956: d <= 8'h00; 15'h6957: d <= 8'h00;
                15'h6958: d <= 8'h45; 15'h6959: d <= 8'h35; 15'h695A: d <= 8'h32; 15'h695B: d <= 8'h00;
                15'h695C: d <= 8'h00; 15'h695D: d <= 8'h00; 15'h695E: d <= 8'h00; 15'h695F: d <= 8'h00;
                15'h6960: d <= 8'h00; 15'h6961: d <= 8'h00; 15'h6962: d <= 8'h00; 15'h6963: d <= 8'h00;
                15'h6964: d <= 8'h00; 15'h6965: d <= 8'h00; 15'h6966: d <= 8'h00; 15'h6967: d <= 8'h00;
                15'h6968: d <= 8'h00; 15'h6969: d <= 8'h00; 15'h696A: d <= 8'h00; 15'h696B: d <= 8'h00;
                15'h696C: d <= 8'h00; 15'h696D: d <= 8'h00; 15'h696E: d <= 8'h00; 15'h696F: d <= 8'h00;
                15'h6970: d <= 8'h00; 15'h6971: d <= 8'h00; 15'h6972: d <= 8'h00; 15'h6973: d <= 8'h00;
                15'h6974: d <= 8'h00; 15'h6975: d <= 8'h00; 15'h6976: d <= 8'h00; 15'h6977: d <= 8'h00;
                15'h6978: d <= 8'h00; 15'h6979: d <= 8'h00; 15'h697A: d <= 8'h00; 15'h697B: d <= 8'h00;
                15'h697C: d <= 8'h00; 15'h697D: d <= 8'h00; 15'h697E: d <= 8'h00; 15'h697F: d <= 8'hE0;
                15'h6980: d <= 8'h10; 15'h6981: d <= 8'h15; 15'h6982: d <= 8'h1A; 15'h6983: d <= 8'h1F;
                15'h6984: d <= 8'h20; 15'h6985: d <= 8'h25; 15'h6986: d <= 8'h2A; 15'h6987: d <= 8'h2F;
                15'h6988: d <= 8'h34; 15'h6989: d <= 8'h38; 15'h698A: d <= 8'h3C; 15'h698B: d <= 8'h31;
                15'h698C: d <= 8'h39; 15'h698D: d <= 8'h3D; 15'h698E: d <= 8'h32; 15'h698F: d <= 8'h36;
                15'h6990: d <= 8'h3E; 15'h6991: d <= 8'h33; 15'h6992: d <= 8'h37; 15'h6993: d <= 8'h3B;
                15'h6994: d <= 8'h44; 15'h6995: d <= 8'h48; 15'h6996: d <= 8'h4C; 15'h6997: d <= 8'h41;
                15'h6998: d <= 8'h49; 15'h6999: d <= 8'h4D; 15'h699A: d <= 8'h42; 15'h699B: d <= 8'h46;
                15'h699C: d <= 8'h4E; 15'h699D: d <= 8'h43; 15'h699E: d <= 8'h47; 15'h699F: d <= 8'h4B;
                15'h69A0: d <= 8'h50; 15'h69A1: d <= 8'h55; 15'h69A2: d <= 8'h5A; 15'h69A3: d <= 8'h5F;
                15'h69A4: d <= 8'h60; 15'h69A5: d <= 8'h65; 15'h69A6: d <= 8'h6A; 15'h69A7: d <= 8'h6F;
                15'h69A8: d <= 8'h74; 15'h69A9: d <= 8'h78; 15'h69AA: d <= 8'h7C; 15'h69AB: d <= 8'h71;
                15'h69AC: d <= 8'h79; 15'h69AD: d <= 8'h7D; 15'h69AE: d <= 8'h72; 15'h69AF: d <= 8'h76;
                15'h69B0: d <= 8'h7E; 15'h69B1: d <= 8'h73; 15'h69B2: d <= 8'h77; 15'h69B3: d <= 8'h7B;
                15'h69B4: d <= 8'h84; 15'h69B5: d <= 8'h88; 15'h69B6: d <= 8'h8C; 15'h69B7: d <= 8'h81;
                15'h69B8: d <= 8'h89; 15'h69B9: d <= 8'h8D; 15'h69BA: d <= 8'h82; 15'h69BB: d <= 8'h86;
                15'h69BC: d <= 8'h8E; 15'h69BD: d <= 8'h83; 15'h69BE: d <= 8'h87; 15'h69BF: d <= 8'h8B;
                15'h69C0: d <= 8'h90; 15'h69C1: d <= 8'h95; 15'h69C2: d <= 8'h9A; 15'h69C3: d <= 8'h9F;
                15'h69C4: d <= 8'hA4; 15'h69C5: d <= 8'hA8; 15'h69C6: d <= 8'hAC; 15'h69C7: d <= 8'hA1;
                15'h69C8: d <= 8'hA9; 15'h69C9: d <= 8'hAD; 15'h69CA: d <= 8'hA2; 15'h69CB: d <= 8'hA6;
                15'h69CC: d <= 8'hAE; 15'h69CD: d <= 8'hA3; 15'h69CE: d <= 8'hA7; 15'h69CF: d <= 8'hAB;
                15'h69D0: d <= 8'hB4; 15'h69D1: d <= 8'hB8; 15'h69D2: d <= 8'hBC; 15'h69D3: d <= 8'hB1;
                15'h69D4: d <= 8'hB9; 15'h69D5: d <= 8'hBD; 15'h69D6: d <= 8'hB2; 15'h69D7: d <= 8'hB6;
                15'h69D8: d <= 8'hBE; 15'h69D9: d <= 8'hB3; 15'h69DA: d <= 8'hB7; 15'h69DB: d <= 8'hBB;
                15'h69DC: d <= 8'hC4; 15'h69DD: d <= 8'hC8; 15'h69DE: d <= 8'hCC; 15'h69DF: d <= 8'hC1;
                15'h69E0: d <= 8'hC9; 15'h69E1: d <= 8'hCD; 15'h69E2: d <= 8'hC2; 15'h69E3: d <= 8'hC6;
                15'h69E4: d <= 8'hCE; 15'h69E5: d <= 8'hC3; 15'h69E6: d <= 8'hC7; 15'h69E7: d <= 8'hCB;
                15'h69E8: d <= 8'hC0; 15'h69E9: d <= 8'hC5; 15'h69EA: d <= 8'hCA; 15'h69EB: d <= 8'hCF;
                15'h69EC: d <= 8'hD0; 15'h69ED: d <= 8'hD5; 15'h69EE: d <= 8'hDA; 15'h69EF: d <= 8'hDF;
                15'h69F0: d <= 8'h74; 15'h69F1: d <= 8'h78; 15'h69F2: d <= 8'h7C; 15'h69F3: d <= 8'h71;
                15'h69F4: d <= 8'h79; 15'h69F5: d <= 8'h7D; 15'h69F6: d <= 8'h72; 15'h69F7: d <= 8'h76;
                15'h69F8: d <= 8'h7E; 15'h69F9: d <= 8'h73; 15'h69FA: d <= 8'h77; 15'h69FB: d <= 8'h7B;
                15'h69FC: d <= 8'hA0; 15'h69FD: d <= 8'hA5; 15'h69FE: d <= 8'hAA; 15'h69FF: d <= 8'hAF;
                15'h6A00: d <= 8'h00; 15'h6A01: d <= 8'h00; 15'h6A02: d <= 8'h00; 15'h6A03: d <= 8'h00;
                15'h6A04: d <= 8'h00; 15'h6A05: d <= 8'h00; 15'h6A06: d <= 8'h00; 15'h6A07: d <= 8'h00;
                15'h6A08: d <= 8'h00; 15'h6A09: d <= 8'h00; 15'h6A0A: d <= 8'h00; 15'h6A0B: d <= 8'h00;
                15'h6A0C: d <= 8'h00; 15'h6A0D: d <= 8'h00; 15'h6A0E: d <= 8'h00; 15'h6A0F: d <= 8'h00;
                15'h6A10: d <= 8'h00; 15'h6A11: d <= 8'h00; 15'h6A12: d <= 8'h00; 15'h6A13: d <= 8'h00;
                15'h6A14: d <= 8'h00; 15'h6A15: d <= 8'h00; 15'h6A16: d <= 8'h00; 15'h6A17: d <= 8'h00;
                15'h6A18: d <= 8'h00; 15'h6A19: d <= 8'h00; 15'h6A1A: d <= 8'h00; 15'h6A1B: d <= 8'h00;
                15'h6A1C: d <= 8'h00; 15'h6A1D: d <= 8'h00; 15'h6A1E: d <= 8'h00; 15'h6A1F: d <= 8'h00;
                15'h6A20: d <= 8'h00; 15'h6A21: d <= 8'h00; 15'h6A22: d <= 8'h00; 15'h6A23: d <= 8'h00;
                15'h6A24: d <= 8'h00; 15'h6A25: d <= 8'h00; 15'h6A26: d <= 8'h00; 15'h6A27: d <= 8'h00;
                15'h6A28: d <= 8'h00; 15'h6A29: d <= 8'h00; 15'h6A2A: d <= 8'h00; 15'h6A2B: d <= 8'h00;
                15'h6A2C: d <= 8'h00; 15'h6A2D: d <= 8'h00; 15'h6A2E: d <= 8'h00; 15'h6A2F: d <= 8'h7B;
                15'h6A30: d <= 8'h00; 15'h6A31: d <= 8'h00; 15'h6A32: d <= 8'h00; 15'h6A33: d <= 8'h00;
                15'h6A34: d <= 8'h00; 15'h6A35: d <= 8'h00; 15'h6A36: d <= 8'h00; 15'h6A37: d <= 8'h00;
                15'h6A38: d <= 8'h00; 15'h6A39: d <= 8'h00; 15'h6A3A: d <= 8'h00; 15'h6A3B: d <= 8'h00;
                15'h6A3C: d <= 8'h00; 15'h6A3D: d <= 8'h00; 15'h6A3E: d <= 8'h00; 15'h6A3F: d <= 8'h00;
                15'h6A40: d <= 8'h00; 15'h6A41: d <= 8'h00; 15'h6A42: d <= 8'h00; 15'h6A43: d <= 8'h00;
                15'h6A44: d <= 8'h00; 15'h6A45: d <= 8'h00; 15'h6A46: d <= 8'h00; 15'h6A47: d <= 8'h00;
                15'h6A48: d <= 8'h00; 15'h6A49: d <= 8'h00; 15'h6A4A: d <= 8'h00; 15'h6A4B: d <= 8'h00;
                15'h6A4C: d <= 8'h00; 15'h6A4D: d <= 8'h00; 15'h6A4E: d <= 8'h00; 15'h6A4F: d <= 8'h00;
                15'h6A50: d <= 8'h00; 15'h6A51: d <= 8'h00; 15'h6A52: d <= 8'h00; 15'h6A53: d <= 8'h00;
                15'h6A54: d <= 8'h00; 15'h6A55: d <= 8'h00; 15'h6A56: d <= 8'h00; 15'h6A57: d <= 8'h00;
                15'h6A58: d <= 8'h45; 15'h6A59: d <= 8'h35; 15'h6A5A: d <= 8'h32; 15'h6A5B: d <= 8'h00;
                15'h6A5C: d <= 8'h00; 15'h6A5D: d <= 8'h00; 15'h6A5E: d <= 8'h00; 15'h6A5F: d <= 8'h00;
                15'h6A60: d <= 8'h00; 15'h6A61: d <= 8'h00; 15'h6A62: d <= 8'h00; 15'h6A63: d <= 8'h00;
                15'h6A64: d <= 8'h00; 15'h6A65: d <= 8'h00; 15'h6A66: d <= 8'h00; 15'h6A67: d <= 8'h00;
                15'h6A68: d <= 8'h00; 15'h6A69: d <= 8'h00; 15'h6A6A: d <= 8'h00; 15'h6A6B: d <= 8'h00;
                15'h6A6C: d <= 8'h00; 15'h6A6D: d <= 8'h00; 15'h6A6E: d <= 8'h00; 15'h6A6F: d <= 8'h00;
                15'h6A70: d <= 8'h00; 15'h6A71: d <= 8'h00; 15'h6A72: d <= 8'h00; 15'h6A73: d <= 8'h00;
                15'h6A74: d <= 8'h00; 15'h6A75: d <= 8'h00; 15'h6A76: d <= 8'h00; 15'h6A77: d <= 8'h00;
                15'h6A78: d <= 8'h00; 15'h6A79: d <= 8'h00; 15'h6A7A: d <= 8'h00; 15'h6A7B: d <= 8'h00;
                15'h6A7C: d <= 8'h00; 15'h6A7D: d <= 8'h00; 15'h6A7E: d <= 8'h00; 15'h6A7F: d <= 8'hE0;
                15'h6A80: d <= 8'h10; 15'h6A81: d <= 8'h15; 15'h6A82: d <= 8'h1A; 15'h6A83: d <= 8'h1F;
                15'h6A84: d <= 8'h20; 15'h6A85: d <= 8'h25; 15'h6A86: d <= 8'h2A; 15'h6A87: d <= 8'h2F;
                15'h6A88: d <= 8'h34; 15'h6A89: d <= 8'h38; 15'h6A8A: d <= 8'h3C; 15'h6A8B: d <= 8'h31;
                15'h6A8C: d <= 8'h39; 15'h6A8D: d <= 8'h3D; 15'h6A8E: d <= 8'h32; 15'h6A8F: d <= 8'h36;
                15'h6A90: d <= 8'h3E; 15'h6A91: d <= 8'h33; 15'h6A92: d <= 8'h37; 15'h6A93: d <= 8'h3B;
                15'h6A94: d <= 8'h44; 15'h6A95: d <= 8'h48; 15'h6A96: d <= 8'h4C; 15'h6A97: d <= 8'h41;
                15'h6A98: d <= 8'h49; 15'h6A99: d <= 8'h4D; 15'h6A9A: d <= 8'h42; 15'h6A9B: d <= 8'h46;
                15'h6A9C: d <= 8'h4E; 15'h6A9D: d <= 8'h43; 15'h6A9E: d <= 8'h47; 15'h6A9F: d <= 8'h4B;
                15'h6AA0: d <= 8'h50; 15'h6AA1: d <= 8'h55; 15'h6AA2: d <= 8'h5A; 15'h6AA3: d <= 8'h5F;
                15'h6AA4: d <= 8'h60; 15'h6AA5: d <= 8'h65; 15'h6AA6: d <= 8'h6A; 15'h6AA7: d <= 8'h6F;
                15'h6AA8: d <= 8'h74; 15'h6AA9: d <= 8'h78; 15'h6AAA: d <= 8'h7C; 15'h6AAB: d <= 8'h71;
                15'h6AAC: d <= 8'h79; 15'h6AAD: d <= 8'h7D; 15'h6AAE: d <= 8'h72; 15'h6AAF: d <= 8'h76;
                15'h6AB0: d <= 8'h7E; 15'h6AB1: d <= 8'h73; 15'h6AB2: d <= 8'h77; 15'h6AB3: d <= 8'h7B;
                15'h6AB4: d <= 8'h84; 15'h6AB5: d <= 8'h88; 15'h6AB6: d <= 8'h8C; 15'h6AB7: d <= 8'h81;
                15'h6AB8: d <= 8'h89; 15'h6AB9: d <= 8'h8D; 15'h6ABA: d <= 8'h82; 15'h6ABB: d <= 8'h86;
                15'h6ABC: d <= 8'h8E; 15'h6ABD: d <= 8'h83; 15'h6ABE: d <= 8'h87; 15'h6ABF: d <= 8'h8B;
                15'h6AC0: d <= 8'h90; 15'h6AC1: d <= 8'h95; 15'h6AC2: d <= 8'h9A; 15'h6AC3: d <= 8'h9F;
                15'h6AC4: d <= 8'hA4; 15'h6AC5: d <= 8'hA8; 15'h6AC6: d <= 8'hAC; 15'h6AC7: d <= 8'hA1;
                15'h6AC8: d <= 8'hA9; 15'h6AC9: d <= 8'hAD; 15'h6ACA: d <= 8'hA2; 15'h6ACB: d <= 8'hA6;
                15'h6ACC: d <= 8'hAE; 15'h6ACD: d <= 8'hA3; 15'h6ACE: d <= 8'hA7; 15'h6ACF: d <= 8'hAB;
                15'h6AD0: d <= 8'hB4; 15'h6AD1: d <= 8'hB8; 15'h6AD2: d <= 8'hBC; 15'h6AD3: d <= 8'hB1;
                15'h6AD4: d <= 8'hB9; 15'h6AD5: d <= 8'hBD; 15'h6AD6: d <= 8'hB2; 15'h6AD7: d <= 8'hB6;
                15'h6AD8: d <= 8'hBE; 15'h6AD9: d <= 8'hB3; 15'h6ADA: d <= 8'hB7; 15'h6ADB: d <= 8'hBB;
                15'h6ADC: d <= 8'hC4; 15'h6ADD: d <= 8'hC8; 15'h6ADE: d <= 8'hCC; 15'h6ADF: d <= 8'hC1;
                15'h6AE0: d <= 8'hC9; 15'h6AE1: d <= 8'hCD; 15'h6AE2: d <= 8'hC2; 15'h6AE3: d <= 8'hC6;
                15'h6AE4: d <= 8'hCE; 15'h6AE5: d <= 8'hC3; 15'h6AE6: d <= 8'hC7; 15'h6AE7: d <= 8'hCB;
                15'h6AE8: d <= 8'hC0; 15'h6AE9: d <= 8'hC5; 15'h6AEA: d <= 8'hCA; 15'h6AEB: d <= 8'hCF;
                15'h6AEC: d <= 8'hD0; 15'h6AED: d <= 8'hD5; 15'h6AEE: d <= 8'hDA; 15'h6AEF: d <= 8'hDF;
                15'h6AF0: d <= 8'h74; 15'h6AF1: d <= 8'h78; 15'h6AF2: d <= 8'h7C; 15'h6AF3: d <= 8'h71;
                15'h6AF4: d <= 8'h79; 15'h6AF5: d <= 8'h7D; 15'h6AF6: d <= 8'h72; 15'h6AF7: d <= 8'h76;
                15'h6AF8: d <= 8'h7E; 15'h6AF9: d <= 8'h73; 15'h6AFA: d <= 8'h77; 15'h6AFB: d <= 8'h7B;
                15'h6AFC: d <= 8'hA0; 15'h6AFD: d <= 8'hA5; 15'h6AFE: d <= 8'hAA; 15'h6AFF: d <= 8'hAF;
                15'h6B00: d <= 8'h00; 15'h6B01: d <= 8'h00; 15'h6B02: d <= 8'h00; 15'h6B03: d <= 8'h00;
                15'h6B04: d <= 8'h00; 15'h6B05: d <= 8'h00; 15'h6B06: d <= 8'h00; 15'h6B07: d <= 8'h00;
                15'h6B08: d <= 8'h00; 15'h6B09: d <= 8'h00; 15'h6B0A: d <= 8'h00; 15'h6B0B: d <= 8'h00;
                15'h6B0C: d <= 8'h00; 15'h6B0D: d <= 8'h00; 15'h6B0E: d <= 8'h00; 15'h6B0F: d <= 8'h00;
                15'h6B10: d <= 8'h00; 15'h6B11: d <= 8'h00; 15'h6B12: d <= 8'h00; 15'h6B13: d <= 8'h00;
                15'h6B14: d <= 8'h00; 15'h6B15: d <= 8'h00; 15'h6B16: d <= 8'h00; 15'h6B17: d <= 8'h00;
                15'h6B18: d <= 8'h00; 15'h6B19: d <= 8'h00; 15'h6B1A: d <= 8'h00; 15'h6B1B: d <= 8'h00;
                15'h6B1C: d <= 8'h00; 15'h6B1D: d <= 8'h00; 15'h6B1E: d <= 8'h00; 15'h6B1F: d <= 8'h00;
                15'h6B20: d <= 8'h00; 15'h6B21: d <= 8'h00; 15'h6B22: d <= 8'h00; 15'h6B23: d <= 8'h00;
                15'h6B24: d <= 8'h00; 15'h6B25: d <= 8'h00; 15'h6B26: d <= 8'h00; 15'h6B27: d <= 8'h00;
                15'h6B28: d <= 8'h00; 15'h6B29: d <= 8'h00; 15'h6B2A: d <= 8'h00; 15'h6B2B: d <= 8'h00;
                15'h6B2C: d <= 8'h00; 15'h6B2D: d <= 8'h00; 15'h6B2E: d <= 8'h00; 15'h6B2F: d <= 8'h7B;
                15'h6B30: d <= 8'h00; 15'h6B31: d <= 8'h00; 15'h6B32: d <= 8'h00; 15'h6B33: d <= 8'h00;
                15'h6B34: d <= 8'h00; 15'h6B35: d <= 8'h00; 15'h6B36: d <= 8'h00; 15'h6B37: d <= 8'h00;
                15'h6B38: d <= 8'h00; 15'h6B39: d <= 8'h00; 15'h6B3A: d <= 8'h00; 15'h6B3B: d <= 8'h00;
                15'h6B3C: d <= 8'h00; 15'h6B3D: d <= 8'h00; 15'h6B3E: d <= 8'h00; 15'h6B3F: d <= 8'h00;
                15'h6B40: d <= 8'h00; 15'h6B41: d <= 8'h00; 15'h6B42: d <= 8'h00; 15'h6B43: d <= 8'h00;
                15'h6B44: d <= 8'h00; 15'h6B45: d <= 8'h00; 15'h6B46: d <= 8'h00; 15'h6B47: d <= 8'h00;
                15'h6B48: d <= 8'h00; 15'h6B49: d <= 8'h00; 15'h6B4A: d <= 8'h00; 15'h6B4B: d <= 8'h00;
                15'h6B4C: d <= 8'h00; 15'h6B4D: d <= 8'h00; 15'h6B4E: d <= 8'h00; 15'h6B4F: d <= 8'h00;
                15'h6B50: d <= 8'h00; 15'h6B51: d <= 8'h00; 15'h6B52: d <= 8'h00; 15'h6B53: d <= 8'h00;
                15'h6B54: d <= 8'h00; 15'h6B55: d <= 8'h00; 15'h6B56: d <= 8'h00; 15'h6B57: d <= 8'h00;
                15'h6B58: d <= 8'h45; 15'h6B59: d <= 8'h35; 15'h6B5A: d <= 8'h32; 15'h6B5B: d <= 8'h00;
                15'h6B5C: d <= 8'h00; 15'h6B5D: d <= 8'h00; 15'h6B5E: d <= 8'h00; 15'h6B5F: d <= 8'h00;
                15'h6B60: d <= 8'h00; 15'h6B61: d <= 8'h00; 15'h6B62: d <= 8'h00; 15'h6B63: d <= 8'h00;
                15'h6B64: d <= 8'h00; 15'h6B65: d <= 8'h00; 15'h6B66: d <= 8'h00; 15'h6B67: d <= 8'h00;
                15'h6B68: d <= 8'h00; 15'h6B69: d <= 8'h00; 15'h6B6A: d <= 8'h00; 15'h6B6B: d <= 8'h00;
                15'h6B6C: d <= 8'h00; 15'h6B6D: d <= 8'h00; 15'h6B6E: d <= 8'h00; 15'h6B6F: d <= 8'h00;
                15'h6B70: d <= 8'h00; 15'h6B71: d <= 8'h00; 15'h6B72: d <= 8'h00; 15'h6B73: d <= 8'h00;
                15'h6B74: d <= 8'h00; 15'h6B75: d <= 8'h00; 15'h6B76: d <= 8'h00; 15'h6B77: d <= 8'h00;
                15'h6B78: d <= 8'h00; 15'h6B79: d <= 8'h00; 15'h6B7A: d <= 8'h00; 15'h6B7B: d <= 8'h00;
                15'h6B7C: d <= 8'h00; 15'h6B7D: d <= 8'h00; 15'h6B7E: d <= 8'h00; 15'h6B7F: d <= 8'hE0;
                15'h6B80: d <= 8'h10; 15'h6B81: d <= 8'h15; 15'h6B82: d <= 8'h1A; 15'h6B83: d <= 8'h1F;
                15'h6B84: d <= 8'h20; 15'h6B85: d <= 8'h25; 15'h6B86: d <= 8'h2A; 15'h6B87: d <= 8'h2F;
                15'h6B88: d <= 8'h34; 15'h6B89: d <= 8'h38; 15'h6B8A: d <= 8'h3C; 15'h6B8B: d <= 8'h31;
                15'h6B8C: d <= 8'h39; 15'h6B8D: d <= 8'h3D; 15'h6B8E: d <= 8'h32; 15'h6B8F: d <= 8'h36;
                15'h6B90: d <= 8'h3E; 15'h6B91: d <= 8'h33; 15'h6B92: d <= 8'h37; 15'h6B93: d <= 8'h3B;
                15'h6B94: d <= 8'h44; 15'h6B95: d <= 8'h48; 15'h6B96: d <= 8'h4C; 15'h6B97: d <= 8'h41;
                15'h6B98: d <= 8'h49; 15'h6B99: d <= 8'h4D; 15'h6B9A: d <= 8'h42; 15'h6B9B: d <= 8'h46;
                15'h6B9C: d <= 8'h4E; 15'h6B9D: d <= 8'h43; 15'h6B9E: d <= 8'h47; 15'h6B9F: d <= 8'h4B;
                15'h6BA0: d <= 8'h50; 15'h6BA1: d <= 8'h55; 15'h6BA2: d <= 8'h5A; 15'h6BA3: d <= 8'h5F;
                15'h6BA4: d <= 8'h60; 15'h6BA5: d <= 8'h65; 15'h6BA6: d <= 8'h6A; 15'h6BA7: d <= 8'h6F;
                15'h6BA8: d <= 8'h74; 15'h6BA9: d <= 8'h78; 15'h6BAA: d <= 8'h7C; 15'h6BAB: d <= 8'h71;
                15'h6BAC: d <= 8'h79; 15'h6BAD: d <= 8'h7D; 15'h6BAE: d <= 8'h72; 15'h6BAF: d <= 8'h76;
                15'h6BB0: d <= 8'h7E; 15'h6BB1: d <= 8'h73; 15'h6BB2: d <= 8'h77; 15'h6BB3: d <= 8'h7B;
                15'h6BB4: d <= 8'h84; 15'h6BB5: d <= 8'h88; 15'h6BB6: d <= 8'h8C; 15'h6BB7: d <= 8'h81;
                15'h6BB8: d <= 8'h89; 15'h6BB9: d <= 8'h8D; 15'h6BBA: d <= 8'h82; 15'h6BBB: d <= 8'h86;
                15'h6BBC: d <= 8'h8E; 15'h6BBD: d <= 8'h83; 15'h6BBE: d <= 8'h87; 15'h6BBF: d <= 8'h8B;
                15'h6BC0: d <= 8'h90; 15'h6BC1: d <= 8'h95; 15'h6BC2: d <= 8'h9A; 15'h6BC3: d <= 8'h9F;
                15'h6BC4: d <= 8'hA4; 15'h6BC5: d <= 8'hA8; 15'h6BC6: d <= 8'hAC; 15'h6BC7: d <= 8'hA1;
                15'h6BC8: d <= 8'hA9; 15'h6BC9: d <= 8'hAD; 15'h6BCA: d <= 8'hA2; 15'h6BCB: d <= 8'hA6;
                15'h6BCC: d <= 8'hAE; 15'h6BCD: d <= 8'hA3; 15'h6BCE: d <= 8'hA7; 15'h6BCF: d <= 8'hAB;
                15'h6BD0: d <= 8'hB4; 15'h6BD1: d <= 8'hB8; 15'h6BD2: d <= 8'hBC; 15'h6BD3: d <= 8'hB1;
                15'h6BD4: d <= 8'hB9; 15'h6BD5: d <= 8'hBD; 15'h6BD6: d <= 8'hB2; 15'h6BD7: d <= 8'hB6;
                15'h6BD8: d <= 8'hBE; 15'h6BD9: d <= 8'hB3; 15'h6BDA: d <= 8'hB7; 15'h6BDB: d <= 8'hBB;
                15'h6BDC: d <= 8'hC4; 15'h6BDD: d <= 8'hC8; 15'h6BDE: d <= 8'hCC; 15'h6BDF: d <= 8'hC1;
                15'h6BE0: d <= 8'hC9; 15'h6BE1: d <= 8'hCD; 15'h6BE2: d <= 8'hC2; 15'h6BE3: d <= 8'hC6;
                15'h6BE4: d <= 8'hCE; 15'h6BE5: d <= 8'hC3; 15'h6BE6: d <= 8'hC7; 15'h6BE7: d <= 8'hCB;
                15'h6BE8: d <= 8'hC0; 15'h6BE9: d <= 8'hC5; 15'h6BEA: d <= 8'hCA; 15'h6BEB: d <= 8'hCF;
                15'h6BEC: d <= 8'hD0; 15'h6BED: d <= 8'hD5; 15'h6BEE: d <= 8'hDA; 15'h6BEF: d <= 8'hDF;
                15'h6BF0: d <= 8'h74; 15'h6BF1: d <= 8'h78; 15'h6BF2: d <= 8'h7C; 15'h6BF3: d <= 8'h71;
                15'h6BF4: d <= 8'h79; 15'h6BF5: d <= 8'h7D; 15'h6BF6: d <= 8'h72; 15'h6BF7: d <= 8'h76;
                15'h6BF8: d <= 8'h7E; 15'h6BF9: d <= 8'h73; 15'h6BFA: d <= 8'h77; 15'h6BFB: d <= 8'h7B;
                15'h6BFC: d <= 8'hA0; 15'h6BFD: d <= 8'hA5; 15'h6BFE: d <= 8'hAA; 15'h6BFF: d <= 8'hAF;
                15'h6C00: d <= 8'h00; 15'h6C01: d <= 8'h00; 15'h6C02: d <= 8'h00; 15'h6C03: d <= 8'h00;
                15'h6C04: d <= 8'h00; 15'h6C05: d <= 8'h00; 15'h6C06: d <= 8'h00; 15'h6C07: d <= 8'h00;
                15'h6C08: d <= 8'h00; 15'h6C09: d <= 8'h00; 15'h6C0A: d <= 8'h00; 15'h6C0B: d <= 8'h00;
                15'h6C0C: d <= 8'h00; 15'h6C0D: d <= 8'h00; 15'h6C0E: d <= 8'h00; 15'h6C0F: d <= 8'h00;
                15'h6C10: d <= 8'h00; 15'h6C11: d <= 8'h00; 15'h6C12: d <= 8'h00; 15'h6C13: d <= 8'h00;
                15'h6C14: d <= 8'h00; 15'h6C15: d <= 8'h00; 15'h6C16: d <= 8'h00; 15'h6C17: d <= 8'h00;
                15'h6C18: d <= 8'h00; 15'h6C19: d <= 8'h00; 15'h6C1A: d <= 8'h00; 15'h6C1B: d <= 8'h00;
                15'h6C1C: d <= 8'h00; 15'h6C1D: d <= 8'h00; 15'h6C1E: d <= 8'h00; 15'h6C1F: d <= 8'h00;
                15'h6C20: d <= 8'h00; 15'h6C21: d <= 8'h00; 15'h6C22: d <= 8'h00; 15'h6C23: d <= 8'h00;
                15'h6C24: d <= 8'h00; 15'h6C25: d <= 8'h00; 15'h6C26: d <= 8'h00; 15'h6C27: d <= 8'h00;
                15'h6C28: d <= 8'h00; 15'h6C29: d <= 8'h00; 15'h6C2A: d <= 8'h00; 15'h6C2B: d <= 8'h00;
                15'h6C2C: d <= 8'h00; 15'h6C2D: d <= 8'h00; 15'h6C2E: d <= 8'h00; 15'h6C2F: d <= 8'h7B;
                15'h6C30: d <= 8'h00; 15'h6C31: d <= 8'h00; 15'h6C32: d <= 8'h00; 15'h6C33: d <= 8'h00;
                15'h6C34: d <= 8'h00; 15'h6C35: d <= 8'h00; 15'h6C36: d <= 8'h00; 15'h6C37: d <= 8'h00;
                15'h6C38: d <= 8'h00; 15'h6C39: d <= 8'h00; 15'h6C3A: d <= 8'h00; 15'h6C3B: d <= 8'h00;
                15'h6C3C: d <= 8'h00; 15'h6C3D: d <= 8'h00; 15'h6C3E: d <= 8'h00; 15'h6C3F: d <= 8'h00;
                15'h6C40: d <= 8'h00; 15'h6C41: d <= 8'h00; 15'h6C42: d <= 8'h00; 15'h6C43: d <= 8'h00;
                15'h6C44: d <= 8'h00; 15'h6C45: d <= 8'h00; 15'h6C46: d <= 8'h00; 15'h6C47: d <= 8'h00;
                15'h6C48: d <= 8'h00; 15'h6C49: d <= 8'h00; 15'h6C4A: d <= 8'h00; 15'h6C4B: d <= 8'h00;
                15'h6C4C: d <= 8'h00; 15'h6C4D: d <= 8'h00; 15'h6C4E: d <= 8'h00; 15'h6C4F: d <= 8'h00;
                15'h6C50: d <= 8'h00; 15'h6C51: d <= 8'h00; 15'h6C52: d <= 8'h00; 15'h6C53: d <= 8'h00;
                15'h6C54: d <= 8'h00; 15'h6C55: d <= 8'h00; 15'h6C56: d <= 8'h00; 15'h6C57: d <= 8'h00;
                15'h6C58: d <= 8'h45; 15'h6C59: d <= 8'h35; 15'h6C5A: d <= 8'h32; 15'h6C5B: d <= 8'h00;
                15'h6C5C: d <= 8'h00; 15'h6C5D: d <= 8'h00; 15'h6C5E: d <= 8'h00; 15'h6C5F: d <= 8'h00;
                15'h6C60: d <= 8'h00; 15'h6C61: d <= 8'h00; 15'h6C62: d <= 8'h00; 15'h6C63: d <= 8'h00;
                15'h6C64: d <= 8'h00; 15'h6C65: d <= 8'h00; 15'h6C66: d <= 8'h00; 15'h6C67: d <= 8'h00;
                15'h6C68: d <= 8'h00; 15'h6C69: d <= 8'h00; 15'h6C6A: d <= 8'h00; 15'h6C6B: d <= 8'h00;
                15'h6C6C: d <= 8'h00; 15'h6C6D: d <= 8'h00; 15'h6C6E: d <= 8'h00; 15'h6C6F: d <= 8'h00;
                15'h6C70: d <= 8'h00; 15'h6C71: d <= 8'h00; 15'h6C72: d <= 8'h00; 15'h6C73: d <= 8'h00;
                15'h6C74: d <= 8'h00; 15'h6C75: d <= 8'h00; 15'h6C76: d <= 8'h00; 15'h6C77: d <= 8'h00;
                15'h6C78: d <= 8'h00; 15'h6C79: d <= 8'h00; 15'h6C7A: d <= 8'h00; 15'h6C7B: d <= 8'h00;
                15'h6C7C: d <= 8'h00; 15'h6C7D: d <= 8'h00; 15'h6C7E: d <= 8'h00; 15'h6C7F: d <= 8'hE0;
                15'h6C80: d <= 8'h10; 15'h6C81: d <= 8'h15; 15'h6C82: d <= 8'h1A; 15'h6C83: d <= 8'h1F;
                15'h6C84: d <= 8'h20; 15'h6C85: d <= 8'h25; 15'h6C86: d <= 8'h2A; 15'h6C87: d <= 8'h2F;
                15'h6C88: d <= 8'h34; 15'h6C89: d <= 8'h38; 15'h6C8A: d <= 8'h3C; 15'h6C8B: d <= 8'h31;
                15'h6C8C: d <= 8'h39; 15'h6C8D: d <= 8'h3D; 15'h6C8E: d <= 8'h32; 15'h6C8F: d <= 8'h36;
                15'h6C90: d <= 8'h3E; 15'h6C91: d <= 8'h33; 15'h6C92: d <= 8'h37; 15'h6C93: d <= 8'h3B;
                15'h6C94: d <= 8'h44; 15'h6C95: d <= 8'h48; 15'h6C96: d <= 8'h4C; 15'h6C97: d <= 8'h41;
                15'h6C98: d <= 8'h49; 15'h6C99: d <= 8'h4D; 15'h6C9A: d <= 8'h42; 15'h6C9B: d <= 8'h46;
                15'h6C9C: d <= 8'h4E; 15'h6C9D: d <= 8'h43; 15'h6C9E: d <= 8'h47; 15'h6C9F: d <= 8'h4B;
                15'h6CA0: d <= 8'h50; 15'h6CA1: d <= 8'h55; 15'h6CA2: d <= 8'h5A; 15'h6CA3: d <= 8'h5F;
                15'h6CA4: d <= 8'h60; 15'h6CA5: d <= 8'h65; 15'h6CA6: d <= 8'h6A; 15'h6CA7: d <= 8'h6F;
                15'h6CA8: d <= 8'h74; 15'h6CA9: d <= 8'h78; 15'h6CAA: d <= 8'h7C; 15'h6CAB: d <= 8'h71;
                15'h6CAC: d <= 8'h79; 15'h6CAD: d <= 8'h7D; 15'h6CAE: d <= 8'h72; 15'h6CAF: d <= 8'h76;
                15'h6CB0: d <= 8'h7E; 15'h6CB1: d <= 8'h73; 15'h6CB2: d <= 8'h77; 15'h6CB3: d <= 8'h7B;
                15'h6CB4: d <= 8'h84; 15'h6CB5: d <= 8'h88; 15'h6CB6: d <= 8'h8C; 15'h6CB7: d <= 8'h81;
                15'h6CB8: d <= 8'h89; 15'h6CB9: d <= 8'h8D; 15'h6CBA: d <= 8'h82; 15'h6CBB: d <= 8'h86;
                15'h6CBC: d <= 8'h8E; 15'h6CBD: d <= 8'h83; 15'h6CBE: d <= 8'h87; 15'h6CBF: d <= 8'h8B;
                15'h6CC0: d <= 8'h90; 15'h6CC1: d <= 8'h95; 15'h6CC2: d <= 8'h9A; 15'h6CC3: d <= 8'h9F;
                15'h6CC4: d <= 8'hA4; 15'h6CC5: d <= 8'hA8; 15'h6CC6: d <= 8'hAC; 15'h6CC7: d <= 8'hA1;
                15'h6CC8: d <= 8'hA9; 15'h6CC9: d <= 8'hAD; 15'h6CCA: d <= 8'hA2; 15'h6CCB: d <= 8'hA6;
                15'h6CCC: d <= 8'hAE; 15'h6CCD: d <= 8'hA3; 15'h6CCE: d <= 8'hA7; 15'h6CCF: d <= 8'hAB;
                15'h6CD0: d <= 8'hB4; 15'h6CD1: d <= 8'hB8; 15'h6CD2: d <= 8'hBC; 15'h6CD3: d <= 8'hB1;
                15'h6CD4: d <= 8'hB9; 15'h6CD5: d <= 8'hBD; 15'h6CD6: d <= 8'hB2; 15'h6CD7: d <= 8'hB6;
                15'h6CD8: d <= 8'hBE; 15'h6CD9: d <= 8'hB3; 15'h6CDA: d <= 8'hB7; 15'h6CDB: d <= 8'hBB;
                15'h6CDC: d <= 8'hC4; 15'h6CDD: d <= 8'hC8; 15'h6CDE: d <= 8'hCC; 15'h6CDF: d <= 8'hC1;
                15'h6CE0: d <= 8'hC9; 15'h6CE1: d <= 8'hCD; 15'h6CE2: d <= 8'hC2; 15'h6CE3: d <= 8'hC6;
                15'h6CE4: d <= 8'hCE; 15'h6CE5: d <= 8'hC3; 15'h6CE6: d <= 8'hC7; 15'h6CE7: d <= 8'hCB;
                15'h6CE8: d <= 8'hC0; 15'h6CE9: d <= 8'hC5; 15'h6CEA: d <= 8'hCA; 15'h6CEB: d <= 8'hCF;
                15'h6CEC: d <= 8'hD0; 15'h6CED: d <= 8'hD5; 15'h6CEE: d <= 8'hDA; 15'h6CEF: d <= 8'hDF;
                15'h6CF0: d <= 8'h74; 15'h6CF1: d <= 8'h78; 15'h6CF2: d <= 8'h7C; 15'h6CF3: d <= 8'h71;
                15'h6CF4: d <= 8'h79; 15'h6CF5: d <= 8'h7D; 15'h6CF6: d <= 8'h72; 15'h6CF7: d <= 8'h76;
                15'h6CF8: d <= 8'h7E; 15'h6CF9: d <= 8'h73; 15'h6CFA: d <= 8'h77; 15'h6CFB: d <= 8'h7B;
                15'h6CFC: d <= 8'hA0; 15'h6CFD: d <= 8'hA5; 15'h6CFE: d <= 8'hAA; 15'h6CFF: d <= 8'hAF;
                15'h6D00: d <= 8'h00; 15'h6D01: d <= 8'h00; 15'h6D02: d <= 8'h00; 15'h6D03: d <= 8'h00;
                15'h6D04: d <= 8'h00; 15'h6D05: d <= 8'h00; 15'h6D06: d <= 8'h00; 15'h6D07: d <= 8'h00;
                15'h6D08: d <= 8'h00; 15'h6D09: d <= 8'h00; 15'h6D0A: d <= 8'h00; 15'h6D0B: d <= 8'h00;
                15'h6D0C: d <= 8'h00; 15'h6D0D: d <= 8'h00; 15'h6D0E: d <= 8'h00; 15'h6D0F: d <= 8'h00;
                15'h6D10: d <= 8'h00; 15'h6D11: d <= 8'h00; 15'h6D12: d <= 8'h00; 15'h6D13: d <= 8'h00;
                15'h6D14: d <= 8'h00; 15'h6D15: d <= 8'h00; 15'h6D16: d <= 8'h00; 15'h6D17: d <= 8'h00;
                15'h6D18: d <= 8'h00; 15'h6D19: d <= 8'h00; 15'h6D1A: d <= 8'h00; 15'h6D1B: d <= 8'h00;
                15'h6D1C: d <= 8'h00; 15'h6D1D: d <= 8'h00; 15'h6D1E: d <= 8'h00; 15'h6D1F: d <= 8'h00;
                15'h6D20: d <= 8'h00; 15'h6D21: d <= 8'h00; 15'h6D22: d <= 8'h00; 15'h6D23: d <= 8'h00;
                15'h6D24: d <= 8'h00; 15'h6D25: d <= 8'h00; 15'h6D26: d <= 8'h00; 15'h6D27: d <= 8'h00;
                15'h6D28: d <= 8'h00; 15'h6D29: d <= 8'h00; 15'h6D2A: d <= 8'h00; 15'h6D2B: d <= 8'h00;
                15'h6D2C: d <= 8'h00; 15'h6D2D: d <= 8'h00; 15'h6D2E: d <= 8'h00; 15'h6D2F: d <= 8'h7B;
                15'h6D30: d <= 8'h00; 15'h6D31: d <= 8'h00; 15'h6D32: d <= 8'h00; 15'h6D33: d <= 8'h00;
                15'h6D34: d <= 8'h00; 15'h6D35: d <= 8'h00; 15'h6D36: d <= 8'h00; 15'h6D37: d <= 8'h00;
                15'h6D38: d <= 8'h00; 15'h6D39: d <= 8'h00; 15'h6D3A: d <= 8'h00; 15'h6D3B: d <= 8'h00;
                15'h6D3C: d <= 8'h00; 15'h6D3D: d <= 8'h00; 15'h6D3E: d <= 8'h00; 15'h6D3F: d <= 8'h00;
                15'h6D40: d <= 8'h00; 15'h6D41: d <= 8'h00; 15'h6D42: d <= 8'h00; 15'h6D43: d <= 8'h00;
                15'h6D44: d <= 8'h00; 15'h6D45: d <= 8'h00; 15'h6D46: d <= 8'h00; 15'h6D47: d <= 8'h00;
                15'h6D48: d <= 8'h00; 15'h6D49: d <= 8'h00; 15'h6D4A: d <= 8'h00; 15'h6D4B: d <= 8'h00;
                15'h6D4C: d <= 8'h00; 15'h6D4D: d <= 8'h00; 15'h6D4E: d <= 8'h00; 15'h6D4F: d <= 8'h00;
                15'h6D50: d <= 8'h00; 15'h6D51: d <= 8'h00; 15'h6D52: d <= 8'h00; 15'h6D53: d <= 8'h00;
                15'h6D54: d <= 8'h00; 15'h6D55: d <= 8'h00; 15'h6D56: d <= 8'h00; 15'h6D57: d <= 8'h00;
                15'h6D58: d <= 8'h45; 15'h6D59: d <= 8'h35; 15'h6D5A: d <= 8'h32; 15'h6D5B: d <= 8'h00;
                15'h6D5C: d <= 8'h00; 15'h6D5D: d <= 8'h00; 15'h6D5E: d <= 8'h00; 15'h6D5F: d <= 8'h00;
                15'h6D60: d <= 8'h00; 15'h6D61: d <= 8'h00; 15'h6D62: d <= 8'h00; 15'h6D63: d <= 8'h00;
                15'h6D64: d <= 8'h00; 15'h6D65: d <= 8'h00; 15'h6D66: d <= 8'h00; 15'h6D67: d <= 8'h00;
                15'h6D68: d <= 8'h00; 15'h6D69: d <= 8'h00; 15'h6D6A: d <= 8'h00; 15'h6D6B: d <= 8'h00;
                15'h6D6C: d <= 8'h00; 15'h6D6D: d <= 8'h00; 15'h6D6E: d <= 8'h00; 15'h6D6F: d <= 8'h00;
                15'h6D70: d <= 8'h00; 15'h6D71: d <= 8'h00; 15'h6D72: d <= 8'h00; 15'h6D73: d <= 8'h00;
                15'h6D74: d <= 8'h00; 15'h6D75: d <= 8'h00; 15'h6D76: d <= 8'h00; 15'h6D77: d <= 8'h00;
                15'h6D78: d <= 8'h00; 15'h6D79: d <= 8'h00; 15'h6D7A: d <= 8'h00; 15'h6D7B: d <= 8'h00;
                15'h6D7C: d <= 8'h00; 15'h6D7D: d <= 8'h00; 15'h6D7E: d <= 8'h00; 15'h6D7F: d <= 8'hE0;
                15'h6D80: d <= 8'h10; 15'h6D81: d <= 8'h15; 15'h6D82: d <= 8'h1A; 15'h6D83: d <= 8'h1F;
                15'h6D84: d <= 8'h20; 15'h6D85: d <= 8'h25; 15'h6D86: d <= 8'h2A; 15'h6D87: d <= 8'h2F;
                15'h6D88: d <= 8'h34; 15'h6D89: d <= 8'h38; 15'h6D8A: d <= 8'h3C; 15'h6D8B: d <= 8'h31;
                15'h6D8C: d <= 8'h39; 15'h6D8D: d <= 8'h3D; 15'h6D8E: d <= 8'h32; 15'h6D8F: d <= 8'h36;
                15'h6D90: d <= 8'h3E; 15'h6D91: d <= 8'h33; 15'h6D92: d <= 8'h37; 15'h6D93: d <= 8'h3B;
                15'h6D94: d <= 8'h44; 15'h6D95: d <= 8'h48; 15'h6D96: d <= 8'h4C; 15'h6D97: d <= 8'h41;
                15'h6D98: d <= 8'h49; 15'h6D99: d <= 8'h4D; 15'h6D9A: d <= 8'h42; 15'h6D9B: d <= 8'h46;
                15'h6D9C: d <= 8'h4E; 15'h6D9D: d <= 8'h43; 15'h6D9E: d <= 8'h47; 15'h6D9F: d <= 8'h4B;
                15'h6DA0: d <= 8'h50; 15'h6DA1: d <= 8'h55; 15'h6DA2: d <= 8'h5A; 15'h6DA3: d <= 8'h5F;
                15'h6DA4: d <= 8'h60; 15'h6DA5: d <= 8'h65; 15'h6DA6: d <= 8'h6A; 15'h6DA7: d <= 8'h6F;
                15'h6DA8: d <= 8'h74; 15'h6DA9: d <= 8'h78; 15'h6DAA: d <= 8'h7C; 15'h6DAB: d <= 8'h71;
                15'h6DAC: d <= 8'h79; 15'h6DAD: d <= 8'h7D; 15'h6DAE: d <= 8'h72; 15'h6DAF: d <= 8'h76;
                15'h6DB0: d <= 8'h7E; 15'h6DB1: d <= 8'h73; 15'h6DB2: d <= 8'h77; 15'h6DB3: d <= 8'h7B;
                15'h6DB4: d <= 8'h84; 15'h6DB5: d <= 8'h88; 15'h6DB6: d <= 8'h8C; 15'h6DB7: d <= 8'h81;
                15'h6DB8: d <= 8'h89; 15'h6DB9: d <= 8'h8D; 15'h6DBA: d <= 8'h82; 15'h6DBB: d <= 8'h86;
                15'h6DBC: d <= 8'h8E; 15'h6DBD: d <= 8'h83; 15'h6DBE: d <= 8'h87; 15'h6DBF: d <= 8'h8B;
                15'h6DC0: d <= 8'h90; 15'h6DC1: d <= 8'h95; 15'h6DC2: d <= 8'h9A; 15'h6DC3: d <= 8'h9F;
                15'h6DC4: d <= 8'hA4; 15'h6DC5: d <= 8'hA8; 15'h6DC6: d <= 8'hAC; 15'h6DC7: d <= 8'hA1;
                15'h6DC8: d <= 8'hA9; 15'h6DC9: d <= 8'hAD; 15'h6DCA: d <= 8'hA2; 15'h6DCB: d <= 8'hA6;
                15'h6DCC: d <= 8'hAE; 15'h6DCD: d <= 8'hA3; 15'h6DCE: d <= 8'hA7; 15'h6DCF: d <= 8'hAB;
                15'h6DD0: d <= 8'hB4; 15'h6DD1: d <= 8'hB8; 15'h6DD2: d <= 8'hBC; 15'h6DD3: d <= 8'hB1;
                15'h6DD4: d <= 8'hB9; 15'h6DD5: d <= 8'hBD; 15'h6DD6: d <= 8'hB2; 15'h6DD7: d <= 8'hB6;
                15'h6DD8: d <= 8'hBE; 15'h6DD9: d <= 8'hB3; 15'h6DDA: d <= 8'hB7; 15'h6DDB: d <= 8'hBB;
                15'h6DDC: d <= 8'hC4; 15'h6DDD: d <= 8'hC8; 15'h6DDE: d <= 8'hCC; 15'h6DDF: d <= 8'hC1;
                15'h6DE0: d <= 8'hC9; 15'h6DE1: d <= 8'hCD; 15'h6DE2: d <= 8'hC2; 15'h6DE3: d <= 8'hC6;
                15'h6DE4: d <= 8'hCE; 15'h6DE5: d <= 8'hC3; 15'h6DE6: d <= 8'hC7; 15'h6DE7: d <= 8'hCB;
                15'h6DE8: d <= 8'hC0; 15'h6DE9: d <= 8'hC5; 15'h6DEA: d <= 8'hCA; 15'h6DEB: d <= 8'hCF;
                15'h6DEC: d <= 8'hD0; 15'h6DED: d <= 8'hD5; 15'h6DEE: d <= 8'hDA; 15'h6DEF: d <= 8'hDF;
                15'h6DF0: d <= 8'h74; 15'h6DF1: d <= 8'h78; 15'h6DF2: d <= 8'h7C; 15'h6DF3: d <= 8'h71;
                15'h6DF4: d <= 8'h79; 15'h6DF5: d <= 8'h7D; 15'h6DF6: d <= 8'h72; 15'h6DF7: d <= 8'h76;
                15'h6DF8: d <= 8'h7E; 15'h6DF9: d <= 8'h73; 15'h6DFA: d <= 8'h77; 15'h6DFB: d <= 8'h7B;
                15'h6DFC: d <= 8'hA0; 15'h6DFD: d <= 8'hA5; 15'h6DFE: d <= 8'hAA; 15'h6DFF: d <= 8'hAF;
                15'h6E00: d <= 8'h00; 15'h6E01: d <= 8'h00; 15'h6E02: d <= 8'h00; 15'h6E03: d <= 8'h00;
                15'h6E04: d <= 8'h00; 15'h6E05: d <= 8'h00; 15'h6E06: d <= 8'h00; 15'h6E07: d <= 8'h00;
                15'h6E08: d <= 8'h00; 15'h6E09: d <= 8'h00; 15'h6E0A: d <= 8'h00; 15'h6E0B: d <= 8'h00;
                15'h6E0C: d <= 8'h00; 15'h6E0D: d <= 8'h00; 15'h6E0E: d <= 8'h00; 15'h6E0F: d <= 8'h00;
                15'h6E10: d <= 8'h00; 15'h6E11: d <= 8'h00; 15'h6E12: d <= 8'h00; 15'h6E13: d <= 8'h00;
                15'h6E14: d <= 8'h00; 15'h6E15: d <= 8'h00; 15'h6E16: d <= 8'h00; 15'h6E17: d <= 8'h00;
                15'h6E18: d <= 8'h00; 15'h6E19: d <= 8'h00; 15'h6E1A: d <= 8'h00; 15'h6E1B: d <= 8'h00;
                15'h6E1C: d <= 8'h00; 15'h6E1D: d <= 8'h00; 15'h6E1E: d <= 8'h00; 15'h6E1F: d <= 8'h00;
                15'h6E20: d <= 8'h00; 15'h6E21: d <= 8'h00; 15'h6E22: d <= 8'h00; 15'h6E23: d <= 8'h00;
                15'h6E24: d <= 8'h00; 15'h6E25: d <= 8'h00; 15'h6E26: d <= 8'h00; 15'h6E27: d <= 8'h00;
                15'h6E28: d <= 8'h00; 15'h6E29: d <= 8'h00; 15'h6E2A: d <= 8'h00; 15'h6E2B: d <= 8'h00;
                15'h6E2C: d <= 8'h00; 15'h6E2D: d <= 8'h00; 15'h6E2E: d <= 8'h00; 15'h6E2F: d <= 8'h7B;
                15'h6E30: d <= 8'h00; 15'h6E31: d <= 8'h00; 15'h6E32: d <= 8'h00; 15'h6E33: d <= 8'h00;
                15'h6E34: d <= 8'h00; 15'h6E35: d <= 8'h00; 15'h6E36: d <= 8'h00; 15'h6E37: d <= 8'h00;
                15'h6E38: d <= 8'h00; 15'h6E39: d <= 8'h00; 15'h6E3A: d <= 8'h00; 15'h6E3B: d <= 8'h00;
                15'h6E3C: d <= 8'h00; 15'h6E3D: d <= 8'h00; 15'h6E3E: d <= 8'h00; 15'h6E3F: d <= 8'h00;
                15'h6E40: d <= 8'h00; 15'h6E41: d <= 8'h00; 15'h6E42: d <= 8'h00; 15'h6E43: d <= 8'h00;
                15'h6E44: d <= 8'h00; 15'h6E45: d <= 8'h00; 15'h6E46: d <= 8'h00; 15'h6E47: d <= 8'h00;
                15'h6E48: d <= 8'h00; 15'h6E49: d <= 8'h00; 15'h6E4A: d <= 8'h00; 15'h6E4B: d <= 8'h00;
                15'h6E4C: d <= 8'h00; 15'h6E4D: d <= 8'h00; 15'h6E4E: d <= 8'h00; 15'h6E4F: d <= 8'h00;
                15'h6E50: d <= 8'h00; 15'h6E51: d <= 8'h00; 15'h6E52: d <= 8'h00; 15'h6E53: d <= 8'h00;
                15'h6E54: d <= 8'h00; 15'h6E55: d <= 8'h00; 15'h6E56: d <= 8'h00; 15'h6E57: d <= 8'h00;
                15'h6E58: d <= 8'h45; 15'h6E59: d <= 8'h35; 15'h6E5A: d <= 8'h32; 15'h6E5B: d <= 8'h00;
                15'h6E5C: d <= 8'h00; 15'h6E5D: d <= 8'h00; 15'h6E5E: d <= 8'h00; 15'h6E5F: d <= 8'h00;
                15'h6E60: d <= 8'h00; 15'h6E61: d <= 8'h00; 15'h6E62: d <= 8'h00; 15'h6E63: d <= 8'h00;
                15'h6E64: d <= 8'h00; 15'h6E65: d <= 8'h00; 15'h6E66: d <= 8'h00; 15'h6E67: d <= 8'h00;
                15'h6E68: d <= 8'h00; 15'h6E69: d <= 8'h00; 15'h6E6A: d <= 8'h00; 15'h6E6B: d <= 8'h00;
                15'h6E6C: d <= 8'h00; 15'h6E6D: d <= 8'h00; 15'h6E6E: d <= 8'h00; 15'h6E6F: d <= 8'h00;
                15'h6E70: d <= 8'h00; 15'h6E71: d <= 8'h00; 15'h6E72: d <= 8'h00; 15'h6E73: d <= 8'h00;
                15'h6E74: d <= 8'h00; 15'h6E75: d <= 8'h00; 15'h6E76: d <= 8'h00; 15'h6E77: d <= 8'h00;
                15'h6E78: d <= 8'h00; 15'h6E79: d <= 8'h00; 15'h6E7A: d <= 8'h00; 15'h6E7B: d <= 8'h00;
                15'h6E7C: d <= 8'h00; 15'h6E7D: d <= 8'h00; 15'h6E7E: d <= 8'h00; 15'h6E7F: d <= 8'hE0;
                15'h6E80: d <= 8'h10; 15'h6E81: d <= 8'h15; 15'h6E82: d <= 8'h1A; 15'h6E83: d <= 8'h1F;
                15'h6E84: d <= 8'h20; 15'h6E85: d <= 8'h25; 15'h6E86: d <= 8'h2A; 15'h6E87: d <= 8'h2F;
                15'h6E88: d <= 8'h34; 15'h6E89: d <= 8'h38; 15'h6E8A: d <= 8'h3C; 15'h6E8B: d <= 8'h31;
                15'h6E8C: d <= 8'h39; 15'h6E8D: d <= 8'h3D; 15'h6E8E: d <= 8'h32; 15'h6E8F: d <= 8'h36;
                15'h6E90: d <= 8'h3E; 15'h6E91: d <= 8'h33; 15'h6E92: d <= 8'h37; 15'h6E93: d <= 8'h3B;
                15'h6E94: d <= 8'h44; 15'h6E95: d <= 8'h48; 15'h6E96: d <= 8'h4C; 15'h6E97: d <= 8'h41;
                15'h6E98: d <= 8'h49; 15'h6E99: d <= 8'h4D; 15'h6E9A: d <= 8'h42; 15'h6E9B: d <= 8'h46;
                15'h6E9C: d <= 8'h4E; 15'h6E9D: d <= 8'h43; 15'h6E9E: d <= 8'h47; 15'h6E9F: d <= 8'h4B;
                15'h6EA0: d <= 8'h50; 15'h6EA1: d <= 8'h55; 15'h6EA2: d <= 8'h5A; 15'h6EA3: d <= 8'h5F;
                15'h6EA4: d <= 8'h60; 15'h6EA5: d <= 8'h65; 15'h6EA6: d <= 8'h6A; 15'h6EA7: d <= 8'h6F;
                15'h6EA8: d <= 8'h74; 15'h6EA9: d <= 8'h78; 15'h6EAA: d <= 8'h7C; 15'h6EAB: d <= 8'h71;
                15'h6EAC: d <= 8'h79; 15'h6EAD: d <= 8'h7D; 15'h6EAE: d <= 8'h72; 15'h6EAF: d <= 8'h76;
                15'h6EB0: d <= 8'h7E; 15'h6EB1: d <= 8'h73; 15'h6EB2: d <= 8'h77; 15'h6EB3: d <= 8'h7B;
                15'h6EB4: d <= 8'h84; 15'h6EB5: d <= 8'h88; 15'h6EB6: d <= 8'h8C; 15'h6EB7: d <= 8'h81;
                15'h6EB8: d <= 8'h89; 15'h6EB9: d <= 8'h8D; 15'h6EBA: d <= 8'h82; 15'h6EBB: d <= 8'h86;
                15'h6EBC: d <= 8'h8E; 15'h6EBD: d <= 8'h83; 15'h6EBE: d <= 8'h87; 15'h6EBF: d <= 8'h8B;
                15'h6EC0: d <= 8'h90; 15'h6EC1: d <= 8'h95; 15'h6EC2: d <= 8'h9A; 15'h6EC3: d <= 8'h9F;
                15'h6EC4: d <= 8'hA4; 15'h6EC5: d <= 8'hA8; 15'h6EC6: d <= 8'hAC; 15'h6EC7: d <= 8'hA1;
                15'h6EC8: d <= 8'hA9; 15'h6EC9: d <= 8'hAD; 15'h6ECA: d <= 8'hA2; 15'h6ECB: d <= 8'hA6;
                15'h6ECC: d <= 8'hAE; 15'h6ECD: d <= 8'hA3; 15'h6ECE: d <= 8'hA7; 15'h6ECF: d <= 8'hAB;
                15'h6ED0: d <= 8'hB4; 15'h6ED1: d <= 8'hB8; 15'h6ED2: d <= 8'hBC; 15'h6ED3: d <= 8'hB1;
                15'h6ED4: d <= 8'hB9; 15'h6ED5: d <= 8'hBD; 15'h6ED6: d <= 8'hB2; 15'h6ED7: d <= 8'hB6;
                15'h6ED8: d <= 8'hBE; 15'h6ED9: d <= 8'hB3; 15'h6EDA: d <= 8'hB7; 15'h6EDB: d <= 8'hBB;
                15'h6EDC: d <= 8'hC4; 15'h6EDD: d <= 8'hC8; 15'h6EDE: d <= 8'hCC; 15'h6EDF: d <= 8'hC1;
                15'h6EE0: d <= 8'hC9; 15'h6EE1: d <= 8'hCD; 15'h6EE2: d <= 8'hC2; 15'h6EE3: d <= 8'hC6;
                15'h6EE4: d <= 8'hCE; 15'h6EE5: d <= 8'hC3; 15'h6EE6: d <= 8'hC7; 15'h6EE7: d <= 8'hCB;
                15'h6EE8: d <= 8'hC0; 15'h6EE9: d <= 8'hC5; 15'h6EEA: d <= 8'hCA; 15'h6EEB: d <= 8'hCF;
                15'h6EEC: d <= 8'hD0; 15'h6EED: d <= 8'hD5; 15'h6EEE: d <= 8'hDA; 15'h6EEF: d <= 8'hDF;
                15'h6EF0: d <= 8'h74; 15'h6EF1: d <= 8'h78; 15'h6EF2: d <= 8'h7C; 15'h6EF3: d <= 8'h71;
                15'h6EF4: d <= 8'h79; 15'h6EF5: d <= 8'h7D; 15'h6EF6: d <= 8'h72; 15'h6EF7: d <= 8'h76;
                15'h6EF8: d <= 8'h7E; 15'h6EF9: d <= 8'h73; 15'h6EFA: d <= 8'h77; 15'h6EFB: d <= 8'h7B;
                15'h6EFC: d <= 8'hA0; 15'h6EFD: d <= 8'hA5; 15'h6EFE: d <= 8'hAA; 15'h6EFF: d <= 8'hAF;
                15'h6F00: d <= 8'h00; 15'h6F01: d <= 8'h00; 15'h6F02: d <= 8'h00; 15'h6F03: d <= 8'h00;
                15'h6F04: d <= 8'h00; 15'h6F05: d <= 8'h00; 15'h6F06: d <= 8'h00; 15'h6F07: d <= 8'h00;
                15'h6F08: d <= 8'h00; 15'h6F09: d <= 8'h00; 15'h6F0A: d <= 8'h00; 15'h6F0B: d <= 8'h00;
                15'h6F0C: d <= 8'h00; 15'h6F0D: d <= 8'h00; 15'h6F0E: d <= 8'h00; 15'h6F0F: d <= 8'h00;
                15'h6F10: d <= 8'h00; 15'h6F11: d <= 8'h00; 15'h6F12: d <= 8'h00; 15'h6F13: d <= 8'h00;
                15'h6F14: d <= 8'h00; 15'h6F15: d <= 8'h00; 15'h6F16: d <= 8'h00; 15'h6F17: d <= 8'h00;
                15'h6F18: d <= 8'h00; 15'h6F19: d <= 8'h00; 15'h6F1A: d <= 8'h00; 15'h6F1B: d <= 8'h00;
                15'h6F1C: d <= 8'h00; 15'h6F1D: d <= 8'h00; 15'h6F1E: d <= 8'h00; 15'h6F1F: d <= 8'h00;
                15'h6F20: d <= 8'h00; 15'h6F21: d <= 8'h00; 15'h6F22: d <= 8'h00; 15'h6F23: d <= 8'h00;
                15'h6F24: d <= 8'h00; 15'h6F25: d <= 8'h00; 15'h6F26: d <= 8'h00; 15'h6F27: d <= 8'h00;
                15'h6F28: d <= 8'h00; 15'h6F29: d <= 8'h00; 15'h6F2A: d <= 8'h00; 15'h6F2B: d <= 8'h00;
                15'h6F2C: d <= 8'h00; 15'h6F2D: d <= 8'h00; 15'h6F2E: d <= 8'h00; 15'h6F2F: d <= 8'h7B;
                15'h6F30: d <= 8'h00; 15'h6F31: d <= 8'h00; 15'h6F32: d <= 8'h00; 15'h6F33: d <= 8'h00;
                15'h6F34: d <= 8'h00; 15'h6F35: d <= 8'h00; 15'h6F36: d <= 8'h00; 15'h6F37: d <= 8'h00;
                15'h6F38: d <= 8'h00; 15'h6F39: d <= 8'h00; 15'h6F3A: d <= 8'h00; 15'h6F3B: d <= 8'h00;
                15'h6F3C: d <= 8'h00; 15'h6F3D: d <= 8'h00; 15'h6F3E: d <= 8'h00; 15'h6F3F: d <= 8'h00;
                15'h6F40: d <= 8'h00; 15'h6F41: d <= 8'h00; 15'h6F42: d <= 8'h00; 15'h6F43: d <= 8'h00;
                15'h6F44: d <= 8'h00; 15'h6F45: d <= 8'h00; 15'h6F46: d <= 8'h00; 15'h6F47: d <= 8'h00;
                15'h6F48: d <= 8'h00; 15'h6F49: d <= 8'h00; 15'h6F4A: d <= 8'h00; 15'h6F4B: d <= 8'h00;
                15'h6F4C: d <= 8'h00; 15'h6F4D: d <= 8'h00; 15'h6F4E: d <= 8'h00; 15'h6F4F: d <= 8'h00;
                15'h6F50: d <= 8'h00; 15'h6F51: d <= 8'h00; 15'h6F52: d <= 8'h00; 15'h6F53: d <= 8'h00;
                15'h6F54: d <= 8'h00; 15'h6F55: d <= 8'h00; 15'h6F56: d <= 8'h00; 15'h6F57: d <= 8'h00;
                15'h6F58: d <= 8'h45; 15'h6F59: d <= 8'h35; 15'h6F5A: d <= 8'h32; 15'h6F5B: d <= 8'h00;
                15'h6F5C: d <= 8'h00; 15'h6F5D: d <= 8'h00; 15'h6F5E: d <= 8'h00; 15'h6F5F: d <= 8'h00;
                15'h6F60: d <= 8'h00; 15'h6F61: d <= 8'h00; 15'h6F62: d <= 8'h00; 15'h6F63: d <= 8'h00;
                15'h6F64: d <= 8'h00; 15'h6F65: d <= 8'h00; 15'h6F66: d <= 8'h00; 15'h6F67: d <= 8'h00;
                15'h6F68: d <= 8'h00; 15'h6F69: d <= 8'h00; 15'h6F6A: d <= 8'h00; 15'h6F6B: d <= 8'h00;
                15'h6F6C: d <= 8'h00; 15'h6F6D: d <= 8'h00; 15'h6F6E: d <= 8'h00; 15'h6F6F: d <= 8'h00;
                15'h6F70: d <= 8'h00; 15'h6F71: d <= 8'h00; 15'h6F72: d <= 8'h00; 15'h6F73: d <= 8'h00;
                15'h6F74: d <= 8'h00; 15'h6F75: d <= 8'h00; 15'h6F76: d <= 8'h00; 15'h6F77: d <= 8'h00;
                15'h6F78: d <= 8'h00; 15'h6F79: d <= 8'h00; 15'h6F7A: d <= 8'h00; 15'h6F7B: d <= 8'h00;
                15'h6F7C: d <= 8'h00; 15'h6F7D: d <= 8'h00; 15'h6F7E: d <= 8'h00; 15'h6F7F: d <= 8'hE0;
                15'h6F80: d <= 8'h10; 15'h6F81: d <= 8'h15; 15'h6F82: d <= 8'h1A; 15'h6F83: d <= 8'h1F;
                15'h6F84: d <= 8'h20; 15'h6F85: d <= 8'h25; 15'h6F86: d <= 8'h2A; 15'h6F87: d <= 8'h2F;
                15'h6F88: d <= 8'h34; 15'h6F89: d <= 8'h38; 15'h6F8A: d <= 8'h3C; 15'h6F8B: d <= 8'h31;
                15'h6F8C: d <= 8'h39; 15'h6F8D: d <= 8'h3D; 15'h6F8E: d <= 8'h32; 15'h6F8F: d <= 8'h36;
                15'h6F90: d <= 8'h3E; 15'h6F91: d <= 8'h33; 15'h6F92: d <= 8'h37; 15'h6F93: d <= 8'h3B;
                15'h6F94: d <= 8'h44; 15'h6F95: d <= 8'h48; 15'h6F96: d <= 8'h4C; 15'h6F97: d <= 8'h41;
                15'h6F98: d <= 8'h49; 15'h6F99: d <= 8'h4D; 15'h6F9A: d <= 8'h42; 15'h6F9B: d <= 8'h46;
                15'h6F9C: d <= 8'h4E; 15'h6F9D: d <= 8'h43; 15'h6F9E: d <= 8'h47; 15'h6F9F: d <= 8'h4B;
                15'h6FA0: d <= 8'h50; 15'h6FA1: d <= 8'h55; 15'h6FA2: d <= 8'h5A; 15'h6FA3: d <= 8'h5F;
                15'h6FA4: d <= 8'h60; 15'h6FA5: d <= 8'h65; 15'h6FA6: d <= 8'h6A; 15'h6FA7: d <= 8'h6F;
                15'h6FA8: d <= 8'h74; 15'h6FA9: d <= 8'h78; 15'h6FAA: d <= 8'h7C; 15'h6FAB: d <= 8'h71;
                15'h6FAC: d <= 8'h79; 15'h6FAD: d <= 8'h7D; 15'h6FAE: d <= 8'h72; 15'h6FAF: d <= 8'h76;
                15'h6FB0: d <= 8'h7E; 15'h6FB1: d <= 8'h73; 15'h6FB2: d <= 8'h77; 15'h6FB3: d <= 8'h7B;
                15'h6FB4: d <= 8'h84; 15'h6FB5: d <= 8'h88; 15'h6FB6: d <= 8'h8C; 15'h6FB7: d <= 8'h81;
                15'h6FB8: d <= 8'h89; 15'h6FB9: d <= 8'h8D; 15'h6FBA: d <= 8'h82; 15'h6FBB: d <= 8'h86;
                15'h6FBC: d <= 8'h8E; 15'h6FBD: d <= 8'h83; 15'h6FBE: d <= 8'h87; 15'h6FBF: d <= 8'h8B;
                15'h6FC0: d <= 8'h90; 15'h6FC1: d <= 8'h95; 15'h6FC2: d <= 8'h9A; 15'h6FC3: d <= 8'h9F;
                15'h6FC4: d <= 8'hA4; 15'h6FC5: d <= 8'hA8; 15'h6FC6: d <= 8'hAC; 15'h6FC7: d <= 8'hA1;
                15'h6FC8: d <= 8'hA9; 15'h6FC9: d <= 8'hAD; 15'h6FCA: d <= 8'hA2; 15'h6FCB: d <= 8'hA6;
                15'h6FCC: d <= 8'hAE; 15'h6FCD: d <= 8'hA3; 15'h6FCE: d <= 8'hA7; 15'h6FCF: d <= 8'hAB;
                15'h6FD0: d <= 8'hB4; 15'h6FD1: d <= 8'hB8; 15'h6FD2: d <= 8'hBC; 15'h6FD3: d <= 8'hB1;
                15'h6FD4: d <= 8'hB9; 15'h6FD5: d <= 8'hBD; 15'h6FD6: d <= 8'hB2; 15'h6FD7: d <= 8'hB6;
                15'h6FD8: d <= 8'hBE; 15'h6FD9: d <= 8'hB3; 15'h6FDA: d <= 8'hB7; 15'h6FDB: d <= 8'hBB;
                15'h6FDC: d <= 8'hC4; 15'h6FDD: d <= 8'hC8; 15'h6FDE: d <= 8'hCC; 15'h6FDF: d <= 8'hC1;
                15'h6FE0: d <= 8'hC9; 15'h6FE1: d <= 8'hCD; 15'h6FE2: d <= 8'hC2; 15'h6FE3: d <= 8'hC6;
                15'h6FE4: d <= 8'hCE; 15'h6FE5: d <= 8'hC3; 15'h6FE6: d <= 8'hC7; 15'h6FE7: d <= 8'hCB;
                15'h6FE8: d <= 8'hC0; 15'h6FE9: d <= 8'hC5; 15'h6FEA: d <= 8'hCA; 15'h6FEB: d <= 8'hCF;
                15'h6FEC: d <= 8'hD0; 15'h6FED: d <= 8'hD5; 15'h6FEE: d <= 8'hDA; 15'h6FEF: d <= 8'hDF;
                15'h6FF0: d <= 8'h74; 15'h6FF1: d <= 8'h78; 15'h6FF2: d <= 8'h7C; 15'h6FF3: d <= 8'h71;
                15'h6FF4: d <= 8'h79; 15'h6FF5: d <= 8'h7D; 15'h6FF6: d <= 8'h72; 15'h6FF7: d <= 8'h76;
                15'h6FF8: d <= 8'h7E; 15'h6FF9: d <= 8'h73; 15'h6FFA: d <= 8'h77; 15'h6FFB: d <= 8'h7B;
                15'h6FFC: d <= 8'hA0; 15'h6FFD: d <= 8'hA5; 15'h6FFE: d <= 8'hAA; 15'h6FFF: d <= 8'hAF;
                15'h7000: d <= 8'h00; 15'h7001: d <= 8'h00; 15'h7002: d <= 8'h00; 15'h7003: d <= 8'h00;
                15'h7004: d <= 8'h00; 15'h7005: d <= 8'h00; 15'h7006: d <= 8'h00; 15'h7007: d <= 8'h00;
                15'h7008: d <= 8'h00; 15'h7009: d <= 8'h00; 15'h700A: d <= 8'h00; 15'h700B: d <= 8'h00;
                15'h700C: d <= 8'h00; 15'h700D: d <= 8'h00; 15'h700E: d <= 8'h00; 15'h700F: d <= 8'h00;
                15'h7010: d <= 8'h00; 15'h7011: d <= 8'h00; 15'h7012: d <= 8'h00; 15'h7013: d <= 8'h00;
                15'h7014: d <= 8'h00; 15'h7015: d <= 8'h00; 15'h7016: d <= 8'h00; 15'h7017: d <= 8'h00;
                15'h7018: d <= 8'h00; 15'h7019: d <= 8'h00; 15'h701A: d <= 8'h00; 15'h701B: d <= 8'h00;
                15'h701C: d <= 8'h00; 15'h701D: d <= 8'h00; 15'h701E: d <= 8'h00; 15'h701F: d <= 8'h00;
                15'h7020: d <= 8'h00; 15'h7021: d <= 8'h00; 15'h7022: d <= 8'h00; 15'h7023: d <= 8'h00;
                15'h7024: d <= 8'h00; 15'h7025: d <= 8'h00; 15'h7026: d <= 8'h00; 15'h7027: d <= 8'h00;
                15'h7028: d <= 8'h00; 15'h7029: d <= 8'h00; 15'h702A: d <= 8'h00; 15'h702B: d <= 8'h00;
                15'h702C: d <= 8'h00; 15'h702D: d <= 8'h00; 15'h702E: d <= 8'h00; 15'h702F: d <= 8'hAF;
                15'h7030: d <= 8'h00; 15'h7031: d <= 8'h00; 15'h7032: d <= 8'h00; 15'h7033: d <= 8'h00;
                15'h7034: d <= 8'h00; 15'h7035: d <= 8'h00; 15'h7036: d <= 8'h00; 15'h7037: d <= 8'h00;
                15'h7038: d <= 8'h00; 15'h7039: d <= 8'h00; 15'h703A: d <= 8'h00; 15'h703B: d <= 8'h00;
                15'h703C: d <= 8'h00; 15'h703D: d <= 8'h00; 15'h703E: d <= 8'h00; 15'h703F: d <= 8'h00;
                15'h7040: d <= 8'h00; 15'h7041: d <= 8'h00; 15'h7042: d <= 8'h00; 15'h7043: d <= 8'h00;
                15'h7044: d <= 8'h00; 15'h7045: d <= 8'h00; 15'h7046: d <= 8'h00; 15'h7047: d <= 8'h00;
                15'h7048: d <= 8'h00; 15'h7049: d <= 8'h00; 15'h704A: d <= 8'h00; 15'h704B: d <= 8'h00;
                15'h704C: d <= 8'h00; 15'h704D: d <= 8'h00; 15'h704E: d <= 8'h00; 15'h704F: d <= 8'h00;
                15'h7050: d <= 8'h00; 15'h7051: d <= 8'h00; 15'h7052: d <= 8'h00; 15'h7053: d <= 8'h00;
                15'h7054: d <= 8'h00; 15'h7055: d <= 8'h00; 15'h7056: d <= 8'h00; 15'h7057: d <= 8'h00;
                15'h7058: d <= 8'h45; 15'h7059: d <= 8'h35; 15'h705A: d <= 8'hAA; 15'h705B: d <= 8'h00;
                15'h705C: d <= 8'h00; 15'h705D: d <= 8'h00; 15'h705E: d <= 8'h00; 15'h705F: d <= 8'h00;
                15'h7060: d <= 8'h00; 15'h7061: d <= 8'h00; 15'h7062: d <= 8'h00; 15'h7063: d <= 8'h00;
                15'h7064: d <= 8'h00; 15'h7065: d <= 8'h00; 15'h7066: d <= 8'h00; 15'h7067: d <= 8'h00;
                15'h7068: d <= 8'h00; 15'h7069: d <= 8'h00; 15'h706A: d <= 8'h00; 15'h706B: d <= 8'h00;
                15'h706C: d <= 8'h00; 15'h706D: d <= 8'h00; 15'h706E: d <= 8'h00; 15'h706F: d <= 8'h00;
                15'h7070: d <= 8'h00; 15'h7071: d <= 8'h00; 15'h7072: d <= 8'h00; 15'h7073: d <= 8'h00;
                15'h7074: d <= 8'h00; 15'h7075: d <= 8'h00; 15'h7076: d <= 8'h00; 15'h7077: d <= 8'h00;
                15'h7078: d <= 8'h00; 15'h7079: d <= 8'h00; 15'h707A: d <= 8'h00; 15'h707B: d <= 8'h00;
                15'h707C: d <= 8'h00; 15'h707D: d <= 8'h00; 15'h707E: d <= 8'h00; 15'h707F: d <= 8'hE0;
                15'h7080: d <= 8'h10; 15'h7081: d <= 8'h15; 15'h7082: d <= 8'h1A; 15'h7083: d <= 8'h1F;
                15'h7084: d <= 8'h20; 15'h7085: d <= 8'h25; 15'h7086: d <= 8'h2A; 15'h7087: d <= 8'h2F;
                15'h7088: d <= 8'h34; 15'h7089: d <= 8'h38; 15'h708A: d <= 8'h3C; 15'h708B: d <= 8'h31;
                15'h708C: d <= 8'h39; 15'h708D: d <= 8'h3D; 15'h708E: d <= 8'h32; 15'h708F: d <= 8'h36;
                15'h7090: d <= 8'h3E; 15'h7091: d <= 8'h33; 15'h7092: d <= 8'h37; 15'h7093: d <= 8'h3B;
                15'h7094: d <= 8'h44; 15'h7095: d <= 8'h48; 15'h7096: d <= 8'h4C; 15'h7097: d <= 8'h41;
                15'h7098: d <= 8'h49; 15'h7099: d <= 8'h4D; 15'h709A: d <= 8'h42; 15'h709B: d <= 8'h46;
                15'h709C: d <= 8'h4E; 15'h709D: d <= 8'h43; 15'h709E: d <= 8'h47; 15'h709F: d <= 8'h4B;
                15'h70A0: d <= 8'h50; 15'h70A1: d <= 8'h55; 15'h70A2: d <= 8'h5A; 15'h70A3: d <= 8'h5F;
                15'h70A4: d <= 8'h60; 15'h70A5: d <= 8'h65; 15'h70A6: d <= 8'h6A; 15'h70A7: d <= 8'h6F;
                15'h70A8: d <= 8'h74; 15'h70A9: d <= 8'h78; 15'h70AA: d <= 8'h7C; 15'h70AB: d <= 8'h71;
                15'h70AC: d <= 8'h79; 15'h70AD: d <= 8'h7D; 15'h70AE: d <= 8'h72; 15'h70AF: d <= 8'h76;
                15'h70B0: d <= 8'h7E; 15'h70B1: d <= 8'h73; 15'h70B2: d <= 8'h77; 15'h70B3: d <= 8'h7B;
                15'h70B4: d <= 8'h84; 15'h70B5: d <= 8'h88; 15'h70B6: d <= 8'h8C; 15'h70B7: d <= 8'h81;
                15'h70B8: d <= 8'h89; 15'h70B9: d <= 8'h8D; 15'h70BA: d <= 8'h82; 15'h70BB: d <= 8'h86;
                15'h70BC: d <= 8'h8E; 15'h70BD: d <= 8'h83; 15'h70BE: d <= 8'h87; 15'h70BF: d <= 8'h8B;
                15'h70C0: d <= 8'h90; 15'h70C1: d <= 8'h95; 15'h70C2: d <= 8'h9A; 15'h70C3: d <= 8'h9F;
                15'h70C4: d <= 8'hA4; 15'h70C5: d <= 8'hA8; 15'h70C6: d <= 8'hAC; 15'h70C7: d <= 8'hA1;
                15'h70C8: d <= 8'hA9; 15'h70C9: d <= 8'hAD; 15'h70CA: d <= 8'hA2; 15'h70CB: d <= 8'hA6;
                15'h70CC: d <= 8'hAE; 15'h70CD: d <= 8'hA3; 15'h70CE: d <= 8'hA7; 15'h70CF: d <= 8'hAB;
                15'h70D0: d <= 8'hB4; 15'h70D1: d <= 8'hB8; 15'h70D2: d <= 8'hBC; 15'h70D3: d <= 8'hB1;
                15'h70D4: d <= 8'hB9; 15'h70D5: d <= 8'hBD; 15'h70D6: d <= 8'hB2; 15'h70D7: d <= 8'hB6;
                15'h70D8: d <= 8'hBE; 15'h70D9: d <= 8'hB3; 15'h70DA: d <= 8'hB7; 15'h70DB: d <= 8'hBB;
                15'h70DC: d <= 8'hC4; 15'h70DD: d <= 8'hC8; 15'h70DE: d <= 8'hCC; 15'h70DF: d <= 8'hC1;
                15'h70E0: d <= 8'hC9; 15'h70E1: d <= 8'hCD; 15'h70E2: d <= 8'hC2; 15'h70E3: d <= 8'hC6;
                15'h70E4: d <= 8'hCE; 15'h70E5: d <= 8'hC3; 15'h70E6: d <= 8'hC7; 15'h70E7: d <= 8'hCB;
                15'h70E8: d <= 8'hC0; 15'h70E9: d <= 8'hC5; 15'h70EA: d <= 8'hCA; 15'h70EB: d <= 8'hCF;
                15'h70EC: d <= 8'hD0; 15'h70ED: d <= 8'hD5; 15'h70EE: d <= 8'hDA; 15'h70EF: d <= 8'hDF;
                15'h70F0: d <= 8'h74; 15'h70F1: d <= 8'h78; 15'h70F2: d <= 8'h7C; 15'h70F3: d <= 8'h71;
                15'h70F4: d <= 8'h79; 15'h70F5: d <= 8'h7D; 15'h70F6: d <= 8'h72; 15'h70F7: d <= 8'h76;
                15'h70F8: d <= 8'h7E; 15'h70F9: d <= 8'h73; 15'h70FA: d <= 8'h77; 15'h70FB: d <= 8'h7B;
                15'h70FC: d <= 8'hA0; 15'h70FD: d <= 8'hA5; 15'h70FE: d <= 8'hAA; 15'h70FF: d <= 8'hAF;
                15'h7100: d <= 8'h00; 15'h7101: d <= 8'h00; 15'h7102: d <= 8'h00; 15'h7103: d <= 8'h00;
                15'h7104: d <= 8'h00; 15'h7105: d <= 8'h00; 15'h7106: d <= 8'h00; 15'h7107: d <= 8'h00;
                15'h7108: d <= 8'h00; 15'h7109: d <= 8'h00; 15'h710A: d <= 8'h00; 15'h710B: d <= 8'h00;
                15'h710C: d <= 8'h00; 15'h710D: d <= 8'h00; 15'h710E: d <= 8'h00; 15'h710F: d <= 8'h00;
                15'h7110: d <= 8'h00; 15'h7111: d <= 8'h00; 15'h7112: d <= 8'h00; 15'h7113: d <= 8'h00;
                15'h7114: d <= 8'h00; 15'h7115: d <= 8'h00; 15'h7116: d <= 8'h00; 15'h7117: d <= 8'h00;
                15'h7118: d <= 8'h00; 15'h7119: d <= 8'h00; 15'h711A: d <= 8'h00; 15'h711B: d <= 8'h00;
                15'h711C: d <= 8'h00; 15'h711D: d <= 8'h00; 15'h711E: d <= 8'h00; 15'h711F: d <= 8'h00;
                15'h7120: d <= 8'h00; 15'h7121: d <= 8'h00; 15'h7122: d <= 8'h00; 15'h7123: d <= 8'h00;
                15'h7124: d <= 8'h00; 15'h7125: d <= 8'h00; 15'h7126: d <= 8'h00; 15'h7127: d <= 8'h00;
                15'h7128: d <= 8'h00; 15'h7129: d <= 8'h00; 15'h712A: d <= 8'h00; 15'h712B: d <= 8'h00;
                15'h712C: d <= 8'h00; 15'h712D: d <= 8'h00; 15'h712E: d <= 8'h00; 15'h712F: d <= 8'hAF;
                15'h7130: d <= 8'h00; 15'h7131: d <= 8'h00; 15'h7132: d <= 8'h00; 15'h7133: d <= 8'h00;
                15'h7134: d <= 8'h00; 15'h7135: d <= 8'h00; 15'h7136: d <= 8'h00; 15'h7137: d <= 8'h00;
                15'h7138: d <= 8'h00; 15'h7139: d <= 8'h00; 15'h713A: d <= 8'h00; 15'h713B: d <= 8'h00;
                15'h713C: d <= 8'h00; 15'h713D: d <= 8'h00; 15'h713E: d <= 8'h00; 15'h713F: d <= 8'h00;
                15'h7140: d <= 8'h00; 15'h7141: d <= 8'h00; 15'h7142: d <= 8'h00; 15'h7143: d <= 8'h00;
                15'h7144: d <= 8'h00; 15'h7145: d <= 8'h00; 15'h7146: d <= 8'h00; 15'h7147: d <= 8'h00;
                15'h7148: d <= 8'h00; 15'h7149: d <= 8'h00; 15'h714A: d <= 8'h00; 15'h714B: d <= 8'h00;
                15'h714C: d <= 8'h00; 15'h714D: d <= 8'h00; 15'h714E: d <= 8'h00; 15'h714F: d <= 8'h00;
                15'h7150: d <= 8'h00; 15'h7151: d <= 8'h00; 15'h7152: d <= 8'h00; 15'h7153: d <= 8'h00;
                15'h7154: d <= 8'h00; 15'h7155: d <= 8'h00; 15'h7156: d <= 8'h00; 15'h7157: d <= 8'h00;
                15'h7158: d <= 8'h45; 15'h7159: d <= 8'h35; 15'h715A: d <= 8'hAA; 15'h715B: d <= 8'h00;
                15'h715C: d <= 8'h00; 15'h715D: d <= 8'h00; 15'h715E: d <= 8'h00; 15'h715F: d <= 8'h00;
                15'h7160: d <= 8'h00; 15'h7161: d <= 8'h00; 15'h7162: d <= 8'h00; 15'h7163: d <= 8'h00;
                15'h7164: d <= 8'h00; 15'h7165: d <= 8'h00; 15'h7166: d <= 8'h00; 15'h7167: d <= 8'h00;
                15'h7168: d <= 8'h00; 15'h7169: d <= 8'h00; 15'h716A: d <= 8'h00; 15'h716B: d <= 8'h00;
                15'h716C: d <= 8'h00; 15'h716D: d <= 8'h00; 15'h716E: d <= 8'h00; 15'h716F: d <= 8'h00;
                15'h7170: d <= 8'h00; 15'h7171: d <= 8'h00; 15'h7172: d <= 8'h00; 15'h7173: d <= 8'h00;
                15'h7174: d <= 8'h00; 15'h7175: d <= 8'h00; 15'h7176: d <= 8'h00; 15'h7177: d <= 8'h00;
                15'h7178: d <= 8'h00; 15'h7179: d <= 8'h00; 15'h717A: d <= 8'h00; 15'h717B: d <= 8'h00;
                15'h717C: d <= 8'h00; 15'h717D: d <= 8'h00; 15'h717E: d <= 8'h00; 15'h717F: d <= 8'hE0;
                15'h7180: d <= 8'h10; 15'h7181: d <= 8'h15; 15'h7182: d <= 8'h1A; 15'h7183: d <= 8'h1F;
                15'h7184: d <= 8'h20; 15'h7185: d <= 8'h25; 15'h7186: d <= 8'h2A; 15'h7187: d <= 8'h2F;
                15'h7188: d <= 8'h34; 15'h7189: d <= 8'h38; 15'h718A: d <= 8'h3C; 15'h718B: d <= 8'h31;
                15'h718C: d <= 8'h39; 15'h718D: d <= 8'h3D; 15'h718E: d <= 8'h32; 15'h718F: d <= 8'h36;
                15'h7190: d <= 8'h3E; 15'h7191: d <= 8'h33; 15'h7192: d <= 8'h37; 15'h7193: d <= 8'h3B;
                15'h7194: d <= 8'h44; 15'h7195: d <= 8'h48; 15'h7196: d <= 8'h4C; 15'h7197: d <= 8'h41;
                15'h7198: d <= 8'h49; 15'h7199: d <= 8'h4D; 15'h719A: d <= 8'h42; 15'h719B: d <= 8'h46;
                15'h719C: d <= 8'h4E; 15'h719D: d <= 8'h43; 15'h719E: d <= 8'h47; 15'h719F: d <= 8'h4B;
                15'h71A0: d <= 8'h50; 15'h71A1: d <= 8'h55; 15'h71A2: d <= 8'h5A; 15'h71A3: d <= 8'h5F;
                15'h71A4: d <= 8'h60; 15'h71A5: d <= 8'h65; 15'h71A6: d <= 8'h6A; 15'h71A7: d <= 8'h6F;
                15'h71A8: d <= 8'h74; 15'h71A9: d <= 8'h78; 15'h71AA: d <= 8'h7C; 15'h71AB: d <= 8'h71;
                15'h71AC: d <= 8'h79; 15'h71AD: d <= 8'h7D; 15'h71AE: d <= 8'h72; 15'h71AF: d <= 8'h76;
                15'h71B0: d <= 8'h7E; 15'h71B1: d <= 8'h73; 15'h71B2: d <= 8'h77; 15'h71B3: d <= 8'h7B;
                15'h71B4: d <= 8'h84; 15'h71B5: d <= 8'h88; 15'h71B6: d <= 8'h8C; 15'h71B7: d <= 8'h81;
                15'h71B8: d <= 8'h89; 15'h71B9: d <= 8'h8D; 15'h71BA: d <= 8'h82; 15'h71BB: d <= 8'h86;
                15'h71BC: d <= 8'h8E; 15'h71BD: d <= 8'h83; 15'h71BE: d <= 8'h87; 15'h71BF: d <= 8'h8B;
                15'h71C0: d <= 8'h90; 15'h71C1: d <= 8'h95; 15'h71C2: d <= 8'h9A; 15'h71C3: d <= 8'h9F;
                15'h71C4: d <= 8'hA4; 15'h71C5: d <= 8'hA8; 15'h71C6: d <= 8'hAC; 15'h71C7: d <= 8'hA1;
                15'h71C8: d <= 8'hA9; 15'h71C9: d <= 8'hAD; 15'h71CA: d <= 8'hA2; 15'h71CB: d <= 8'hA6;
                15'h71CC: d <= 8'hAE; 15'h71CD: d <= 8'hA3; 15'h71CE: d <= 8'hA7; 15'h71CF: d <= 8'hAB;
                15'h71D0: d <= 8'hB4; 15'h71D1: d <= 8'hB8; 15'h71D2: d <= 8'hBC; 15'h71D3: d <= 8'hB1;
                15'h71D4: d <= 8'hB9; 15'h71D5: d <= 8'hBD; 15'h71D6: d <= 8'hB2; 15'h71D7: d <= 8'hB6;
                15'h71D8: d <= 8'hBE; 15'h71D9: d <= 8'hB3; 15'h71DA: d <= 8'hB7; 15'h71DB: d <= 8'hBB;
                15'h71DC: d <= 8'hC4; 15'h71DD: d <= 8'hC8; 15'h71DE: d <= 8'hCC; 15'h71DF: d <= 8'hC1;
                15'h71E0: d <= 8'hC9; 15'h71E1: d <= 8'hCD; 15'h71E2: d <= 8'hC2; 15'h71E3: d <= 8'hC6;
                15'h71E4: d <= 8'hCE; 15'h71E5: d <= 8'hC3; 15'h71E6: d <= 8'hC7; 15'h71E7: d <= 8'hCB;
                15'h71E8: d <= 8'hC0; 15'h71E9: d <= 8'hC5; 15'h71EA: d <= 8'hCA; 15'h71EB: d <= 8'hCF;
                15'h71EC: d <= 8'hD0; 15'h71ED: d <= 8'hD5; 15'h71EE: d <= 8'hDA; 15'h71EF: d <= 8'hDF;
                15'h71F0: d <= 8'h74; 15'h71F1: d <= 8'h78; 15'h71F2: d <= 8'h7C; 15'h71F3: d <= 8'h71;
                15'h71F4: d <= 8'h79; 15'h71F5: d <= 8'h7D; 15'h71F6: d <= 8'h72; 15'h71F7: d <= 8'h76;
                15'h71F8: d <= 8'h7E; 15'h71F9: d <= 8'h73; 15'h71FA: d <= 8'h77; 15'h71FB: d <= 8'h7B;
                15'h71FC: d <= 8'hA0; 15'h71FD: d <= 8'hA5; 15'h71FE: d <= 8'hAA; 15'h71FF: d <= 8'hAF;
                15'h7200: d <= 8'h00; 15'h7201: d <= 8'h00; 15'h7202: d <= 8'h00; 15'h7203: d <= 8'h00;
                15'h7204: d <= 8'h00; 15'h7205: d <= 8'h00; 15'h7206: d <= 8'h00; 15'h7207: d <= 8'h00;
                15'h7208: d <= 8'h00; 15'h7209: d <= 8'h00; 15'h720A: d <= 8'h00; 15'h720B: d <= 8'h00;
                15'h720C: d <= 8'h00; 15'h720D: d <= 8'h00; 15'h720E: d <= 8'h00; 15'h720F: d <= 8'h00;
                15'h7210: d <= 8'h00; 15'h7211: d <= 8'h00; 15'h7212: d <= 8'h00; 15'h7213: d <= 8'h00;
                15'h7214: d <= 8'h00; 15'h7215: d <= 8'h00; 15'h7216: d <= 8'h00; 15'h7217: d <= 8'h00;
                15'h7218: d <= 8'h00; 15'h7219: d <= 8'h00; 15'h721A: d <= 8'h00; 15'h721B: d <= 8'h00;
                15'h721C: d <= 8'h00; 15'h721D: d <= 8'h00; 15'h721E: d <= 8'h00; 15'h721F: d <= 8'h00;
                15'h7220: d <= 8'h00; 15'h7221: d <= 8'h00; 15'h7222: d <= 8'h00; 15'h7223: d <= 8'h00;
                15'h7224: d <= 8'h00; 15'h7225: d <= 8'h00; 15'h7226: d <= 8'h00; 15'h7227: d <= 8'h00;
                15'h7228: d <= 8'h00; 15'h7229: d <= 8'h00; 15'h722A: d <= 8'h00; 15'h722B: d <= 8'h00;
                15'h722C: d <= 8'h00; 15'h722D: d <= 8'h00; 15'h722E: d <= 8'h00; 15'h722F: d <= 8'hAF;
                15'h7230: d <= 8'h00; 15'h7231: d <= 8'h00; 15'h7232: d <= 8'h00; 15'h7233: d <= 8'h00;
                15'h7234: d <= 8'h00; 15'h7235: d <= 8'h00; 15'h7236: d <= 8'h00; 15'h7237: d <= 8'h00;
                15'h7238: d <= 8'h00; 15'h7239: d <= 8'h00; 15'h723A: d <= 8'h00; 15'h723B: d <= 8'h00;
                15'h723C: d <= 8'h00; 15'h723D: d <= 8'h00; 15'h723E: d <= 8'h00; 15'h723F: d <= 8'h00;
                15'h7240: d <= 8'h00; 15'h7241: d <= 8'h00; 15'h7242: d <= 8'h00; 15'h7243: d <= 8'h00;
                15'h7244: d <= 8'h00; 15'h7245: d <= 8'h00; 15'h7246: d <= 8'h00; 15'h7247: d <= 8'h00;
                15'h7248: d <= 8'h00; 15'h7249: d <= 8'h00; 15'h724A: d <= 8'h00; 15'h724B: d <= 8'h00;
                15'h724C: d <= 8'h00; 15'h724D: d <= 8'h00; 15'h724E: d <= 8'h00; 15'h724F: d <= 8'h00;
                15'h7250: d <= 8'h00; 15'h7251: d <= 8'h00; 15'h7252: d <= 8'h00; 15'h7253: d <= 8'h00;
                15'h7254: d <= 8'h00; 15'h7255: d <= 8'h00; 15'h7256: d <= 8'h00; 15'h7257: d <= 8'h00;
                15'h7258: d <= 8'h45; 15'h7259: d <= 8'h35; 15'h725A: d <= 8'hAA; 15'h725B: d <= 8'h00;
                15'h725C: d <= 8'h00; 15'h725D: d <= 8'h00; 15'h725E: d <= 8'h00; 15'h725F: d <= 8'h00;
                15'h7260: d <= 8'h00; 15'h7261: d <= 8'h00; 15'h7262: d <= 8'h00; 15'h7263: d <= 8'h00;
                15'h7264: d <= 8'h00; 15'h7265: d <= 8'h00; 15'h7266: d <= 8'h00; 15'h7267: d <= 8'h00;
                15'h7268: d <= 8'h00; 15'h7269: d <= 8'h00; 15'h726A: d <= 8'h00; 15'h726B: d <= 8'h00;
                15'h726C: d <= 8'h00; 15'h726D: d <= 8'h00; 15'h726E: d <= 8'h00; 15'h726F: d <= 8'h00;
                15'h7270: d <= 8'h00; 15'h7271: d <= 8'h00; 15'h7272: d <= 8'h00; 15'h7273: d <= 8'h00;
                15'h7274: d <= 8'h00; 15'h7275: d <= 8'h00; 15'h7276: d <= 8'h00; 15'h7277: d <= 8'h00;
                15'h7278: d <= 8'h00; 15'h7279: d <= 8'h00; 15'h727A: d <= 8'h00; 15'h727B: d <= 8'h00;
                15'h727C: d <= 8'h00; 15'h727D: d <= 8'h00; 15'h727E: d <= 8'h00; 15'h727F: d <= 8'hE0;
                15'h7280: d <= 8'h10; 15'h7281: d <= 8'h15; 15'h7282: d <= 8'h1A; 15'h7283: d <= 8'h1F;
                15'h7284: d <= 8'h20; 15'h7285: d <= 8'h25; 15'h7286: d <= 8'h2A; 15'h7287: d <= 8'h2F;
                15'h7288: d <= 8'h34; 15'h7289: d <= 8'h38; 15'h728A: d <= 8'h3C; 15'h728B: d <= 8'h31;
                15'h728C: d <= 8'h39; 15'h728D: d <= 8'h3D; 15'h728E: d <= 8'h32; 15'h728F: d <= 8'h36;
                15'h7290: d <= 8'h3E; 15'h7291: d <= 8'h33; 15'h7292: d <= 8'h37; 15'h7293: d <= 8'h3B;
                15'h7294: d <= 8'h44; 15'h7295: d <= 8'h48; 15'h7296: d <= 8'h4C; 15'h7297: d <= 8'h41;
                15'h7298: d <= 8'h49; 15'h7299: d <= 8'h4D; 15'h729A: d <= 8'h42; 15'h729B: d <= 8'h46;
                15'h729C: d <= 8'h4E; 15'h729D: d <= 8'h43; 15'h729E: d <= 8'h47; 15'h729F: d <= 8'h4B;
                15'h72A0: d <= 8'h50; 15'h72A1: d <= 8'h55; 15'h72A2: d <= 8'h5A; 15'h72A3: d <= 8'h5F;
                15'h72A4: d <= 8'h60; 15'h72A5: d <= 8'h65; 15'h72A6: d <= 8'h6A; 15'h72A7: d <= 8'h6F;
                15'h72A8: d <= 8'h74; 15'h72A9: d <= 8'h78; 15'h72AA: d <= 8'h7C; 15'h72AB: d <= 8'h71;
                15'h72AC: d <= 8'h79; 15'h72AD: d <= 8'h7D; 15'h72AE: d <= 8'h72; 15'h72AF: d <= 8'h76;
                15'h72B0: d <= 8'h7E; 15'h72B1: d <= 8'h73; 15'h72B2: d <= 8'h77; 15'h72B3: d <= 8'h7B;
                15'h72B4: d <= 8'h84; 15'h72B5: d <= 8'h88; 15'h72B6: d <= 8'h8C; 15'h72B7: d <= 8'h81;
                15'h72B8: d <= 8'h89; 15'h72B9: d <= 8'h8D; 15'h72BA: d <= 8'h82; 15'h72BB: d <= 8'h86;
                15'h72BC: d <= 8'h8E; 15'h72BD: d <= 8'h83; 15'h72BE: d <= 8'h87; 15'h72BF: d <= 8'h8B;
                15'h72C0: d <= 8'h90; 15'h72C1: d <= 8'h95; 15'h72C2: d <= 8'h9A; 15'h72C3: d <= 8'h9F;
                15'h72C4: d <= 8'hA4; 15'h72C5: d <= 8'hA8; 15'h72C6: d <= 8'hAC; 15'h72C7: d <= 8'hA1;
                15'h72C8: d <= 8'hA9; 15'h72C9: d <= 8'hAD; 15'h72CA: d <= 8'hA2; 15'h72CB: d <= 8'hA6;
                15'h72CC: d <= 8'hAE; 15'h72CD: d <= 8'hA3; 15'h72CE: d <= 8'hA7; 15'h72CF: d <= 8'hAB;
                15'h72D0: d <= 8'hB4; 15'h72D1: d <= 8'hB8; 15'h72D2: d <= 8'hBC; 15'h72D3: d <= 8'hB1;
                15'h72D4: d <= 8'hB9; 15'h72D5: d <= 8'hBD; 15'h72D6: d <= 8'hB2; 15'h72D7: d <= 8'hB6;
                15'h72D8: d <= 8'hBE; 15'h72D9: d <= 8'hB3; 15'h72DA: d <= 8'hB7; 15'h72DB: d <= 8'hBB;
                15'h72DC: d <= 8'hC4; 15'h72DD: d <= 8'hC8; 15'h72DE: d <= 8'hCC; 15'h72DF: d <= 8'hC1;
                15'h72E0: d <= 8'hC9; 15'h72E1: d <= 8'hCD; 15'h72E2: d <= 8'hC2; 15'h72E3: d <= 8'hC6;
                15'h72E4: d <= 8'hCE; 15'h72E5: d <= 8'hC3; 15'h72E6: d <= 8'hC7; 15'h72E7: d <= 8'hCB;
                15'h72E8: d <= 8'hC0; 15'h72E9: d <= 8'hC5; 15'h72EA: d <= 8'hCA; 15'h72EB: d <= 8'hCF;
                15'h72EC: d <= 8'hD0; 15'h72ED: d <= 8'hD5; 15'h72EE: d <= 8'hDA; 15'h72EF: d <= 8'hDF;
                15'h72F0: d <= 8'h74; 15'h72F1: d <= 8'h78; 15'h72F2: d <= 8'h7C; 15'h72F3: d <= 8'h71;
                15'h72F4: d <= 8'h79; 15'h72F5: d <= 8'h7D; 15'h72F6: d <= 8'h72; 15'h72F7: d <= 8'h76;
                15'h72F8: d <= 8'h7E; 15'h72F9: d <= 8'h73; 15'h72FA: d <= 8'h77; 15'h72FB: d <= 8'h7B;
                15'h72FC: d <= 8'hA0; 15'h72FD: d <= 8'hA5; 15'h72FE: d <= 8'hAA; 15'h72FF: d <= 8'hAF;
                15'h7300: d <= 8'h00; 15'h7301: d <= 8'h00; 15'h7302: d <= 8'h00; 15'h7303: d <= 8'h00;
                15'h7304: d <= 8'h00; 15'h7305: d <= 8'h00; 15'h7306: d <= 8'h00; 15'h7307: d <= 8'h00;
                15'h7308: d <= 8'h00; 15'h7309: d <= 8'h00; 15'h730A: d <= 8'h00; 15'h730B: d <= 8'h00;
                15'h730C: d <= 8'h00; 15'h730D: d <= 8'h00; 15'h730E: d <= 8'h00; 15'h730F: d <= 8'h00;
                15'h7310: d <= 8'h00; 15'h7311: d <= 8'h00; 15'h7312: d <= 8'h00; 15'h7313: d <= 8'h00;
                15'h7314: d <= 8'h00; 15'h7315: d <= 8'h00; 15'h7316: d <= 8'h00; 15'h7317: d <= 8'h00;
                15'h7318: d <= 8'h00; 15'h7319: d <= 8'h00; 15'h731A: d <= 8'h00; 15'h731B: d <= 8'h00;
                15'h731C: d <= 8'h00; 15'h731D: d <= 8'h00; 15'h731E: d <= 8'h00; 15'h731F: d <= 8'h00;
                15'h7320: d <= 8'h00; 15'h7321: d <= 8'h00; 15'h7322: d <= 8'h00; 15'h7323: d <= 8'h00;
                15'h7324: d <= 8'h00; 15'h7325: d <= 8'h00; 15'h7326: d <= 8'h00; 15'h7327: d <= 8'h00;
                15'h7328: d <= 8'h00; 15'h7329: d <= 8'h00; 15'h732A: d <= 8'h00; 15'h732B: d <= 8'h00;
                15'h732C: d <= 8'h00; 15'h732D: d <= 8'h00; 15'h732E: d <= 8'h00; 15'h732F: d <= 8'hAF;
                15'h7330: d <= 8'h00; 15'h7331: d <= 8'h00; 15'h7332: d <= 8'h00; 15'h7333: d <= 8'h00;
                15'h7334: d <= 8'h00; 15'h7335: d <= 8'h00; 15'h7336: d <= 8'h00; 15'h7337: d <= 8'h00;
                15'h7338: d <= 8'h00; 15'h7339: d <= 8'h00; 15'h733A: d <= 8'h00; 15'h733B: d <= 8'h00;
                15'h733C: d <= 8'h00; 15'h733D: d <= 8'h00; 15'h733E: d <= 8'h00; 15'h733F: d <= 8'h00;
                15'h7340: d <= 8'h00; 15'h7341: d <= 8'h00; 15'h7342: d <= 8'h00; 15'h7343: d <= 8'h00;
                15'h7344: d <= 8'h00; 15'h7345: d <= 8'h00; 15'h7346: d <= 8'h00; 15'h7347: d <= 8'h00;
                15'h7348: d <= 8'h00; 15'h7349: d <= 8'h00; 15'h734A: d <= 8'h00; 15'h734B: d <= 8'h00;
                15'h734C: d <= 8'h00; 15'h734D: d <= 8'h00; 15'h734E: d <= 8'h00; 15'h734F: d <= 8'h00;
                15'h7350: d <= 8'h00; 15'h7351: d <= 8'h00; 15'h7352: d <= 8'h00; 15'h7353: d <= 8'h00;
                15'h7354: d <= 8'h00; 15'h7355: d <= 8'h00; 15'h7356: d <= 8'h00; 15'h7357: d <= 8'h00;
                15'h7358: d <= 8'h45; 15'h7359: d <= 8'h35; 15'h735A: d <= 8'hAA; 15'h735B: d <= 8'h00;
                15'h735C: d <= 8'h00; 15'h735D: d <= 8'h00; 15'h735E: d <= 8'h00; 15'h735F: d <= 8'h00;
                15'h7360: d <= 8'h00; 15'h7361: d <= 8'h00; 15'h7362: d <= 8'h00; 15'h7363: d <= 8'h00;
                15'h7364: d <= 8'h00; 15'h7365: d <= 8'h00; 15'h7366: d <= 8'h00; 15'h7367: d <= 8'h00;
                15'h7368: d <= 8'h00; 15'h7369: d <= 8'h00; 15'h736A: d <= 8'h00; 15'h736B: d <= 8'h00;
                15'h736C: d <= 8'h00; 15'h736D: d <= 8'h00; 15'h736E: d <= 8'h00; 15'h736F: d <= 8'h00;
                15'h7370: d <= 8'h00; 15'h7371: d <= 8'h00; 15'h7372: d <= 8'h00; 15'h7373: d <= 8'h00;
                15'h7374: d <= 8'h00; 15'h7375: d <= 8'h00; 15'h7376: d <= 8'h00; 15'h7377: d <= 8'h00;
                15'h7378: d <= 8'h00; 15'h7379: d <= 8'h00; 15'h737A: d <= 8'h00; 15'h737B: d <= 8'h00;
                15'h737C: d <= 8'h00; 15'h737D: d <= 8'h00; 15'h737E: d <= 8'h00; 15'h737F: d <= 8'hE0;
                15'h7380: d <= 8'h10; 15'h7381: d <= 8'h15; 15'h7382: d <= 8'h1A; 15'h7383: d <= 8'h1F;
                15'h7384: d <= 8'h20; 15'h7385: d <= 8'h25; 15'h7386: d <= 8'h2A; 15'h7387: d <= 8'h2F;
                15'h7388: d <= 8'h34; 15'h7389: d <= 8'h38; 15'h738A: d <= 8'h3C; 15'h738B: d <= 8'h31;
                15'h738C: d <= 8'h39; 15'h738D: d <= 8'h3D; 15'h738E: d <= 8'h32; 15'h738F: d <= 8'h36;
                15'h7390: d <= 8'h3E; 15'h7391: d <= 8'h33; 15'h7392: d <= 8'h37; 15'h7393: d <= 8'h3B;
                15'h7394: d <= 8'h44; 15'h7395: d <= 8'h48; 15'h7396: d <= 8'h4C; 15'h7397: d <= 8'h41;
                15'h7398: d <= 8'h49; 15'h7399: d <= 8'h4D; 15'h739A: d <= 8'h42; 15'h739B: d <= 8'h46;
                15'h739C: d <= 8'h4E; 15'h739D: d <= 8'h43; 15'h739E: d <= 8'h47; 15'h739F: d <= 8'h4B;
                15'h73A0: d <= 8'h50; 15'h73A1: d <= 8'h55; 15'h73A2: d <= 8'h5A; 15'h73A3: d <= 8'h5F;
                15'h73A4: d <= 8'h60; 15'h73A5: d <= 8'h65; 15'h73A6: d <= 8'h6A; 15'h73A7: d <= 8'h6F;
                15'h73A8: d <= 8'h74; 15'h73A9: d <= 8'h78; 15'h73AA: d <= 8'h7C; 15'h73AB: d <= 8'h71;
                15'h73AC: d <= 8'h79; 15'h73AD: d <= 8'h7D; 15'h73AE: d <= 8'h72; 15'h73AF: d <= 8'h76;
                15'h73B0: d <= 8'h7E; 15'h73B1: d <= 8'h73; 15'h73B2: d <= 8'h77; 15'h73B3: d <= 8'h7B;
                15'h73B4: d <= 8'h84; 15'h73B5: d <= 8'h88; 15'h73B6: d <= 8'h8C; 15'h73B7: d <= 8'h81;
                15'h73B8: d <= 8'h89; 15'h73B9: d <= 8'h8D; 15'h73BA: d <= 8'h82; 15'h73BB: d <= 8'h86;
                15'h73BC: d <= 8'h8E; 15'h73BD: d <= 8'h83; 15'h73BE: d <= 8'h87; 15'h73BF: d <= 8'h8B;
                15'h73C0: d <= 8'h90; 15'h73C1: d <= 8'h95; 15'h73C2: d <= 8'h9A; 15'h73C3: d <= 8'h9F;
                15'h73C4: d <= 8'hA4; 15'h73C5: d <= 8'hA8; 15'h73C6: d <= 8'hAC; 15'h73C7: d <= 8'hA1;
                15'h73C8: d <= 8'hA9; 15'h73C9: d <= 8'hAD; 15'h73CA: d <= 8'hA2; 15'h73CB: d <= 8'hA6;
                15'h73CC: d <= 8'hAE; 15'h73CD: d <= 8'hA3; 15'h73CE: d <= 8'hA7; 15'h73CF: d <= 8'hAB;
                15'h73D0: d <= 8'hB4; 15'h73D1: d <= 8'hB8; 15'h73D2: d <= 8'hBC; 15'h73D3: d <= 8'hB1;
                15'h73D4: d <= 8'hB9; 15'h73D5: d <= 8'hBD; 15'h73D6: d <= 8'hB2; 15'h73D7: d <= 8'hB6;
                15'h73D8: d <= 8'hBE; 15'h73D9: d <= 8'hB3; 15'h73DA: d <= 8'hB7; 15'h73DB: d <= 8'hBB;
                15'h73DC: d <= 8'hC4; 15'h73DD: d <= 8'hC8; 15'h73DE: d <= 8'hCC; 15'h73DF: d <= 8'hC1;
                15'h73E0: d <= 8'hC9; 15'h73E1: d <= 8'hCD; 15'h73E2: d <= 8'hC2; 15'h73E3: d <= 8'hC6;
                15'h73E4: d <= 8'hCE; 15'h73E5: d <= 8'hC3; 15'h73E6: d <= 8'hC7; 15'h73E7: d <= 8'hCB;
                15'h73E8: d <= 8'hC0; 15'h73E9: d <= 8'hC5; 15'h73EA: d <= 8'hCA; 15'h73EB: d <= 8'hCF;
                15'h73EC: d <= 8'hD0; 15'h73ED: d <= 8'hD5; 15'h73EE: d <= 8'hDA; 15'h73EF: d <= 8'hDF;
                15'h73F0: d <= 8'h74; 15'h73F1: d <= 8'h78; 15'h73F2: d <= 8'h7C; 15'h73F3: d <= 8'h71;
                15'h73F4: d <= 8'h79; 15'h73F5: d <= 8'h7D; 15'h73F6: d <= 8'h72; 15'h73F7: d <= 8'h76;
                15'h73F8: d <= 8'h7E; 15'h73F9: d <= 8'h73; 15'h73FA: d <= 8'h77; 15'h73FB: d <= 8'h7B;
                15'h73FC: d <= 8'hA0; 15'h73FD: d <= 8'hA5; 15'h73FE: d <= 8'hAA; 15'h73FF: d <= 8'hAF;
                15'h7400: d <= 8'h00; 15'h7401: d <= 8'h00; 15'h7402: d <= 8'h00; 15'h7403: d <= 8'h00;
                15'h7404: d <= 8'h00; 15'h7405: d <= 8'h00; 15'h7406: d <= 8'h00; 15'h7407: d <= 8'h00;
                15'h7408: d <= 8'h00; 15'h7409: d <= 8'h00; 15'h740A: d <= 8'h00; 15'h740B: d <= 8'h00;
                15'h740C: d <= 8'h00; 15'h740D: d <= 8'h00; 15'h740E: d <= 8'h00; 15'h740F: d <= 8'h00;
                15'h7410: d <= 8'h00; 15'h7411: d <= 8'h00; 15'h7412: d <= 8'h00; 15'h7413: d <= 8'h00;
                15'h7414: d <= 8'h00; 15'h7415: d <= 8'h00; 15'h7416: d <= 8'h00; 15'h7417: d <= 8'h00;
                15'h7418: d <= 8'h00; 15'h7419: d <= 8'h00; 15'h741A: d <= 8'h00; 15'h741B: d <= 8'h00;
                15'h741C: d <= 8'h00; 15'h741D: d <= 8'h00; 15'h741E: d <= 8'h00; 15'h741F: d <= 8'h00;
                15'h7420: d <= 8'h00; 15'h7421: d <= 8'h00; 15'h7422: d <= 8'h00; 15'h7423: d <= 8'h00;
                15'h7424: d <= 8'h00; 15'h7425: d <= 8'h00; 15'h7426: d <= 8'h00; 15'h7427: d <= 8'h00;
                15'h7428: d <= 8'h00; 15'h7429: d <= 8'h00; 15'h742A: d <= 8'h00; 15'h742B: d <= 8'h00;
                15'h742C: d <= 8'h00; 15'h742D: d <= 8'h00; 15'h742E: d <= 8'h00; 15'h742F: d <= 8'hAF;
                15'h7430: d <= 8'h00; 15'h7431: d <= 8'h00; 15'h7432: d <= 8'h00; 15'h7433: d <= 8'h00;
                15'h7434: d <= 8'h00; 15'h7435: d <= 8'h00; 15'h7436: d <= 8'h00; 15'h7437: d <= 8'h00;
                15'h7438: d <= 8'h00; 15'h7439: d <= 8'h00; 15'h743A: d <= 8'h00; 15'h743B: d <= 8'h00;
                15'h743C: d <= 8'h00; 15'h743D: d <= 8'h00; 15'h743E: d <= 8'h00; 15'h743F: d <= 8'h00;
                15'h7440: d <= 8'h00; 15'h7441: d <= 8'h00; 15'h7442: d <= 8'h00; 15'h7443: d <= 8'h00;
                15'h7444: d <= 8'h00; 15'h7445: d <= 8'h00; 15'h7446: d <= 8'h00; 15'h7447: d <= 8'h00;
                15'h7448: d <= 8'h00; 15'h7449: d <= 8'h00; 15'h744A: d <= 8'h00; 15'h744B: d <= 8'h00;
                15'h744C: d <= 8'h00; 15'h744D: d <= 8'h00; 15'h744E: d <= 8'h00; 15'h744F: d <= 8'h00;
                15'h7450: d <= 8'h00; 15'h7451: d <= 8'h00; 15'h7452: d <= 8'h00; 15'h7453: d <= 8'h00;
                15'h7454: d <= 8'h00; 15'h7455: d <= 8'h00; 15'h7456: d <= 8'h00; 15'h7457: d <= 8'h00;
                15'h7458: d <= 8'h45; 15'h7459: d <= 8'h35; 15'h745A: d <= 8'hAA; 15'h745B: d <= 8'h00;
                15'h745C: d <= 8'h00; 15'h745D: d <= 8'h00; 15'h745E: d <= 8'h00; 15'h745F: d <= 8'h00;
                15'h7460: d <= 8'h00; 15'h7461: d <= 8'h00; 15'h7462: d <= 8'h00; 15'h7463: d <= 8'h00;
                15'h7464: d <= 8'h00; 15'h7465: d <= 8'h00; 15'h7466: d <= 8'h00; 15'h7467: d <= 8'h00;
                15'h7468: d <= 8'h00; 15'h7469: d <= 8'h00; 15'h746A: d <= 8'h00; 15'h746B: d <= 8'h00;
                15'h746C: d <= 8'h00; 15'h746D: d <= 8'h00; 15'h746E: d <= 8'h00; 15'h746F: d <= 8'h00;
                15'h7470: d <= 8'h00; 15'h7471: d <= 8'h00; 15'h7472: d <= 8'h00; 15'h7473: d <= 8'h00;
                15'h7474: d <= 8'h00; 15'h7475: d <= 8'h00; 15'h7476: d <= 8'h00; 15'h7477: d <= 8'h00;
                15'h7478: d <= 8'h00; 15'h7479: d <= 8'h00; 15'h747A: d <= 8'h00; 15'h747B: d <= 8'h00;
                15'h747C: d <= 8'h00; 15'h747D: d <= 8'h00; 15'h747E: d <= 8'h00; 15'h747F: d <= 8'hE0;
                15'h7480: d <= 8'h10; 15'h7481: d <= 8'h15; 15'h7482: d <= 8'h1A; 15'h7483: d <= 8'h1F;
                15'h7484: d <= 8'h20; 15'h7485: d <= 8'h25; 15'h7486: d <= 8'h2A; 15'h7487: d <= 8'h2F;
                15'h7488: d <= 8'h34; 15'h7489: d <= 8'h38; 15'h748A: d <= 8'h3C; 15'h748B: d <= 8'h31;
                15'h748C: d <= 8'h39; 15'h748D: d <= 8'h3D; 15'h748E: d <= 8'h32; 15'h748F: d <= 8'h36;
                15'h7490: d <= 8'h3E; 15'h7491: d <= 8'h33; 15'h7492: d <= 8'h37; 15'h7493: d <= 8'h3B;
                15'h7494: d <= 8'h44; 15'h7495: d <= 8'h48; 15'h7496: d <= 8'h4C; 15'h7497: d <= 8'h41;
                15'h7498: d <= 8'h49; 15'h7499: d <= 8'h4D; 15'h749A: d <= 8'h42; 15'h749B: d <= 8'h46;
                15'h749C: d <= 8'h4E; 15'h749D: d <= 8'h43; 15'h749E: d <= 8'h47; 15'h749F: d <= 8'h4B;
                15'h74A0: d <= 8'h50; 15'h74A1: d <= 8'h55; 15'h74A2: d <= 8'h5A; 15'h74A3: d <= 8'h5F;
                15'h74A4: d <= 8'h60; 15'h74A5: d <= 8'h65; 15'h74A6: d <= 8'h6A; 15'h74A7: d <= 8'h6F;
                15'h74A8: d <= 8'h74; 15'h74A9: d <= 8'h78; 15'h74AA: d <= 8'h7C; 15'h74AB: d <= 8'h71;
                15'h74AC: d <= 8'h79; 15'h74AD: d <= 8'h7D; 15'h74AE: d <= 8'h72; 15'h74AF: d <= 8'h76;
                15'h74B0: d <= 8'h7E; 15'h74B1: d <= 8'h73; 15'h74B2: d <= 8'h77; 15'h74B3: d <= 8'h7B;
                15'h74B4: d <= 8'h84; 15'h74B5: d <= 8'h88; 15'h74B6: d <= 8'h8C; 15'h74B7: d <= 8'h81;
                15'h74B8: d <= 8'h89; 15'h74B9: d <= 8'h8D; 15'h74BA: d <= 8'h82; 15'h74BB: d <= 8'h86;
                15'h74BC: d <= 8'h8E; 15'h74BD: d <= 8'h83; 15'h74BE: d <= 8'h87; 15'h74BF: d <= 8'h8B;
                15'h74C0: d <= 8'h90; 15'h74C1: d <= 8'h95; 15'h74C2: d <= 8'h9A; 15'h74C3: d <= 8'h9F;
                15'h74C4: d <= 8'hA4; 15'h74C5: d <= 8'hA8; 15'h74C6: d <= 8'hAC; 15'h74C7: d <= 8'hA1;
                15'h74C8: d <= 8'hA9; 15'h74C9: d <= 8'hAD; 15'h74CA: d <= 8'hA2; 15'h74CB: d <= 8'hA6;
                15'h74CC: d <= 8'hAE; 15'h74CD: d <= 8'hA3; 15'h74CE: d <= 8'hA7; 15'h74CF: d <= 8'hAB;
                15'h74D0: d <= 8'hB4; 15'h74D1: d <= 8'hB8; 15'h74D2: d <= 8'hBC; 15'h74D3: d <= 8'hB1;
                15'h74D4: d <= 8'hB9; 15'h74D5: d <= 8'hBD; 15'h74D6: d <= 8'hB2; 15'h74D7: d <= 8'hB6;
                15'h74D8: d <= 8'hBE; 15'h74D9: d <= 8'hB3; 15'h74DA: d <= 8'hB7; 15'h74DB: d <= 8'hBB;
                15'h74DC: d <= 8'hC4; 15'h74DD: d <= 8'hC8; 15'h74DE: d <= 8'hCC; 15'h74DF: d <= 8'hC1;
                15'h74E0: d <= 8'hC9; 15'h74E1: d <= 8'hCD; 15'h74E2: d <= 8'hC2; 15'h74E3: d <= 8'hC6;
                15'h74E4: d <= 8'hCE; 15'h74E5: d <= 8'hC3; 15'h74E6: d <= 8'hC7; 15'h74E7: d <= 8'hCB;
                15'h74E8: d <= 8'hC0; 15'h74E9: d <= 8'hC5; 15'h74EA: d <= 8'hCA; 15'h74EB: d <= 8'hCF;
                15'h74EC: d <= 8'hD0; 15'h74ED: d <= 8'hD5; 15'h74EE: d <= 8'hDA; 15'h74EF: d <= 8'hDF;
                15'h74F0: d <= 8'h74; 15'h74F1: d <= 8'h78; 15'h74F2: d <= 8'h7C; 15'h74F3: d <= 8'h71;
                15'h74F4: d <= 8'h79; 15'h74F5: d <= 8'h7D; 15'h74F6: d <= 8'h72; 15'h74F7: d <= 8'h76;
                15'h74F8: d <= 8'h7E; 15'h74F9: d <= 8'h73; 15'h74FA: d <= 8'h77; 15'h74FB: d <= 8'h7B;
                15'h74FC: d <= 8'hA0; 15'h74FD: d <= 8'hA5; 15'h74FE: d <= 8'hAA; 15'h74FF: d <= 8'hAF;
                15'h7500: d <= 8'h00; 15'h7501: d <= 8'h00; 15'h7502: d <= 8'h00; 15'h7503: d <= 8'h00;
                15'h7504: d <= 8'h00; 15'h7505: d <= 8'h00; 15'h7506: d <= 8'h00; 15'h7507: d <= 8'h00;
                15'h7508: d <= 8'h00; 15'h7509: d <= 8'h00; 15'h750A: d <= 8'h00; 15'h750B: d <= 8'h00;
                15'h750C: d <= 8'h00; 15'h750D: d <= 8'h00; 15'h750E: d <= 8'h00; 15'h750F: d <= 8'h00;
                15'h7510: d <= 8'h00; 15'h7511: d <= 8'h00; 15'h7512: d <= 8'h00; 15'h7513: d <= 8'h00;
                15'h7514: d <= 8'h00; 15'h7515: d <= 8'h00; 15'h7516: d <= 8'h00; 15'h7517: d <= 8'h00;
                15'h7518: d <= 8'h00; 15'h7519: d <= 8'h00; 15'h751A: d <= 8'h00; 15'h751B: d <= 8'h00;
                15'h751C: d <= 8'h00; 15'h751D: d <= 8'h00; 15'h751E: d <= 8'h00; 15'h751F: d <= 8'h00;
                15'h7520: d <= 8'h00; 15'h7521: d <= 8'h00; 15'h7522: d <= 8'h00; 15'h7523: d <= 8'h00;
                15'h7524: d <= 8'h00; 15'h7525: d <= 8'h00; 15'h7526: d <= 8'h00; 15'h7527: d <= 8'h00;
                15'h7528: d <= 8'h00; 15'h7529: d <= 8'h00; 15'h752A: d <= 8'h00; 15'h752B: d <= 8'h00;
                15'h752C: d <= 8'h00; 15'h752D: d <= 8'h00; 15'h752E: d <= 8'h00; 15'h752F: d <= 8'hAF;
                15'h7530: d <= 8'h00; 15'h7531: d <= 8'h00; 15'h7532: d <= 8'h00; 15'h7533: d <= 8'h00;
                15'h7534: d <= 8'h00; 15'h7535: d <= 8'h00; 15'h7536: d <= 8'h00; 15'h7537: d <= 8'h00;
                15'h7538: d <= 8'h00; 15'h7539: d <= 8'h00; 15'h753A: d <= 8'h00; 15'h753B: d <= 8'h00;
                15'h753C: d <= 8'h00; 15'h753D: d <= 8'h00; 15'h753E: d <= 8'h00; 15'h753F: d <= 8'h00;
                15'h7540: d <= 8'h00; 15'h7541: d <= 8'h00; 15'h7542: d <= 8'h00; 15'h7543: d <= 8'h00;
                15'h7544: d <= 8'h00; 15'h7545: d <= 8'h00; 15'h7546: d <= 8'h00; 15'h7547: d <= 8'h00;
                15'h7548: d <= 8'h00; 15'h7549: d <= 8'h00; 15'h754A: d <= 8'h00; 15'h754B: d <= 8'h00;
                15'h754C: d <= 8'h00; 15'h754D: d <= 8'h00; 15'h754E: d <= 8'h00; 15'h754F: d <= 8'h00;
                15'h7550: d <= 8'h00; 15'h7551: d <= 8'h00; 15'h7552: d <= 8'h00; 15'h7553: d <= 8'h00;
                15'h7554: d <= 8'h00; 15'h7555: d <= 8'h00; 15'h7556: d <= 8'h00; 15'h7557: d <= 8'h00;
                15'h7558: d <= 8'h45; 15'h7559: d <= 8'h35; 15'h755A: d <= 8'hAA; 15'h755B: d <= 8'h00;
                15'h755C: d <= 8'h00; 15'h755D: d <= 8'h00; 15'h755E: d <= 8'h00; 15'h755F: d <= 8'h00;
                15'h7560: d <= 8'h00; 15'h7561: d <= 8'h00; 15'h7562: d <= 8'h00; 15'h7563: d <= 8'h00;
                15'h7564: d <= 8'h00; 15'h7565: d <= 8'h00; 15'h7566: d <= 8'h00; 15'h7567: d <= 8'h00;
                15'h7568: d <= 8'h00; 15'h7569: d <= 8'h00; 15'h756A: d <= 8'h00; 15'h756B: d <= 8'h00;
                15'h756C: d <= 8'h00; 15'h756D: d <= 8'h00; 15'h756E: d <= 8'h00; 15'h756F: d <= 8'h00;
                15'h7570: d <= 8'h00; 15'h7571: d <= 8'h00; 15'h7572: d <= 8'h00; 15'h7573: d <= 8'h00;
                15'h7574: d <= 8'h00; 15'h7575: d <= 8'h00; 15'h7576: d <= 8'h00; 15'h7577: d <= 8'h00;
                15'h7578: d <= 8'h00; 15'h7579: d <= 8'h00; 15'h757A: d <= 8'h00; 15'h757B: d <= 8'h00;
                15'h757C: d <= 8'h00; 15'h757D: d <= 8'h00; 15'h757E: d <= 8'h00; 15'h757F: d <= 8'hE0;
                15'h7580: d <= 8'h10; 15'h7581: d <= 8'h15; 15'h7582: d <= 8'h1A; 15'h7583: d <= 8'h1F;
                15'h7584: d <= 8'h20; 15'h7585: d <= 8'h25; 15'h7586: d <= 8'h2A; 15'h7587: d <= 8'h2F;
                15'h7588: d <= 8'h34; 15'h7589: d <= 8'h38; 15'h758A: d <= 8'h3C; 15'h758B: d <= 8'h31;
                15'h758C: d <= 8'h39; 15'h758D: d <= 8'h3D; 15'h758E: d <= 8'h32; 15'h758F: d <= 8'h36;
                15'h7590: d <= 8'h3E; 15'h7591: d <= 8'h33; 15'h7592: d <= 8'h37; 15'h7593: d <= 8'h3B;
                15'h7594: d <= 8'h44; 15'h7595: d <= 8'h48; 15'h7596: d <= 8'h4C; 15'h7597: d <= 8'h41;
                15'h7598: d <= 8'h49; 15'h7599: d <= 8'h4D; 15'h759A: d <= 8'h42; 15'h759B: d <= 8'h46;
                15'h759C: d <= 8'h4E; 15'h759D: d <= 8'h43; 15'h759E: d <= 8'h47; 15'h759F: d <= 8'h4B;
                15'h75A0: d <= 8'h50; 15'h75A1: d <= 8'h55; 15'h75A2: d <= 8'h5A; 15'h75A3: d <= 8'h5F;
                15'h75A4: d <= 8'h60; 15'h75A5: d <= 8'h65; 15'h75A6: d <= 8'h6A; 15'h75A7: d <= 8'h6F;
                15'h75A8: d <= 8'h74; 15'h75A9: d <= 8'h78; 15'h75AA: d <= 8'h7C; 15'h75AB: d <= 8'h71;
                15'h75AC: d <= 8'h79; 15'h75AD: d <= 8'h7D; 15'h75AE: d <= 8'h72; 15'h75AF: d <= 8'h76;
                15'h75B0: d <= 8'h7E; 15'h75B1: d <= 8'h73; 15'h75B2: d <= 8'h77; 15'h75B3: d <= 8'h7B;
                15'h75B4: d <= 8'h84; 15'h75B5: d <= 8'h88; 15'h75B6: d <= 8'h8C; 15'h75B7: d <= 8'h81;
                15'h75B8: d <= 8'h89; 15'h75B9: d <= 8'h8D; 15'h75BA: d <= 8'h82; 15'h75BB: d <= 8'h86;
                15'h75BC: d <= 8'h8E; 15'h75BD: d <= 8'h83; 15'h75BE: d <= 8'h87; 15'h75BF: d <= 8'h8B;
                15'h75C0: d <= 8'h90; 15'h75C1: d <= 8'h95; 15'h75C2: d <= 8'h9A; 15'h75C3: d <= 8'h9F;
                15'h75C4: d <= 8'hA4; 15'h75C5: d <= 8'hA8; 15'h75C6: d <= 8'hAC; 15'h75C7: d <= 8'hA1;
                15'h75C8: d <= 8'hA9; 15'h75C9: d <= 8'hAD; 15'h75CA: d <= 8'hA2; 15'h75CB: d <= 8'hA6;
                15'h75CC: d <= 8'hAE; 15'h75CD: d <= 8'hA3; 15'h75CE: d <= 8'hA7; 15'h75CF: d <= 8'hAB;
                15'h75D0: d <= 8'hB4; 15'h75D1: d <= 8'hB8; 15'h75D2: d <= 8'hBC; 15'h75D3: d <= 8'hB1;
                15'h75D4: d <= 8'hB9; 15'h75D5: d <= 8'hBD; 15'h75D6: d <= 8'hB2; 15'h75D7: d <= 8'hB6;
                15'h75D8: d <= 8'hBE; 15'h75D9: d <= 8'hB3; 15'h75DA: d <= 8'hB7; 15'h75DB: d <= 8'hBB;
                15'h75DC: d <= 8'hC4; 15'h75DD: d <= 8'hC8; 15'h75DE: d <= 8'hCC; 15'h75DF: d <= 8'hC1;
                15'h75E0: d <= 8'hC9; 15'h75E1: d <= 8'hCD; 15'h75E2: d <= 8'hC2; 15'h75E3: d <= 8'hC6;
                15'h75E4: d <= 8'hCE; 15'h75E5: d <= 8'hC3; 15'h75E6: d <= 8'hC7; 15'h75E7: d <= 8'hCB;
                15'h75E8: d <= 8'hC0; 15'h75E9: d <= 8'hC5; 15'h75EA: d <= 8'hCA; 15'h75EB: d <= 8'hCF;
                15'h75EC: d <= 8'hD0; 15'h75ED: d <= 8'hD5; 15'h75EE: d <= 8'hDA; 15'h75EF: d <= 8'hDF;
                15'h75F0: d <= 8'h74; 15'h75F1: d <= 8'h78; 15'h75F2: d <= 8'h7C; 15'h75F3: d <= 8'h71;
                15'h75F4: d <= 8'h79; 15'h75F5: d <= 8'h7D; 15'h75F6: d <= 8'h72; 15'h75F7: d <= 8'h76;
                15'h75F8: d <= 8'h7E; 15'h75F9: d <= 8'h73; 15'h75FA: d <= 8'h77; 15'h75FB: d <= 8'h7B;
                15'h75FC: d <= 8'hA0; 15'h75FD: d <= 8'hA5; 15'h75FE: d <= 8'hAA; 15'h75FF: d <= 8'hAF;
                15'h7600: d <= 8'h00; 15'h7601: d <= 8'h00; 15'h7602: d <= 8'h00; 15'h7603: d <= 8'h00;
                15'h7604: d <= 8'h00; 15'h7605: d <= 8'h00; 15'h7606: d <= 8'h00; 15'h7607: d <= 8'h00;
                15'h7608: d <= 8'h00; 15'h7609: d <= 8'h00; 15'h760A: d <= 8'h00; 15'h760B: d <= 8'h00;
                15'h760C: d <= 8'h00; 15'h760D: d <= 8'h00; 15'h760E: d <= 8'h00; 15'h760F: d <= 8'h00;
                15'h7610: d <= 8'h00; 15'h7611: d <= 8'h00; 15'h7612: d <= 8'h00; 15'h7613: d <= 8'h00;
                15'h7614: d <= 8'h00; 15'h7615: d <= 8'h00; 15'h7616: d <= 8'h00; 15'h7617: d <= 8'h00;
                15'h7618: d <= 8'h00; 15'h7619: d <= 8'h00; 15'h761A: d <= 8'h00; 15'h761B: d <= 8'h00;
                15'h761C: d <= 8'h00; 15'h761D: d <= 8'h00; 15'h761E: d <= 8'h00; 15'h761F: d <= 8'h00;
                15'h7620: d <= 8'h00; 15'h7621: d <= 8'h00; 15'h7622: d <= 8'h00; 15'h7623: d <= 8'h00;
                15'h7624: d <= 8'h00; 15'h7625: d <= 8'h00; 15'h7626: d <= 8'h00; 15'h7627: d <= 8'h00;
                15'h7628: d <= 8'h00; 15'h7629: d <= 8'h00; 15'h762A: d <= 8'h00; 15'h762B: d <= 8'h00;
                15'h762C: d <= 8'h00; 15'h762D: d <= 8'h00; 15'h762E: d <= 8'h00; 15'h762F: d <= 8'hAF;
                15'h7630: d <= 8'h00; 15'h7631: d <= 8'h00; 15'h7632: d <= 8'h00; 15'h7633: d <= 8'h00;
                15'h7634: d <= 8'h00; 15'h7635: d <= 8'h00; 15'h7636: d <= 8'h00; 15'h7637: d <= 8'h00;
                15'h7638: d <= 8'h00; 15'h7639: d <= 8'h00; 15'h763A: d <= 8'h00; 15'h763B: d <= 8'h00;
                15'h763C: d <= 8'h00; 15'h763D: d <= 8'h00; 15'h763E: d <= 8'h00; 15'h763F: d <= 8'h00;
                15'h7640: d <= 8'h00; 15'h7641: d <= 8'h00; 15'h7642: d <= 8'h00; 15'h7643: d <= 8'h00;
                15'h7644: d <= 8'h00; 15'h7645: d <= 8'h00; 15'h7646: d <= 8'h00; 15'h7647: d <= 8'h00;
                15'h7648: d <= 8'h00; 15'h7649: d <= 8'h00; 15'h764A: d <= 8'h00; 15'h764B: d <= 8'h00;
                15'h764C: d <= 8'h00; 15'h764D: d <= 8'h00; 15'h764E: d <= 8'h00; 15'h764F: d <= 8'h00;
                15'h7650: d <= 8'h00; 15'h7651: d <= 8'h00; 15'h7652: d <= 8'h00; 15'h7653: d <= 8'h00;
                15'h7654: d <= 8'h00; 15'h7655: d <= 8'h00; 15'h7656: d <= 8'h00; 15'h7657: d <= 8'h00;
                15'h7658: d <= 8'h45; 15'h7659: d <= 8'h35; 15'h765A: d <= 8'hAA; 15'h765B: d <= 8'h00;
                15'h765C: d <= 8'h00; 15'h765D: d <= 8'h00; 15'h765E: d <= 8'h00; 15'h765F: d <= 8'h00;
                15'h7660: d <= 8'h00; 15'h7661: d <= 8'h00; 15'h7662: d <= 8'h00; 15'h7663: d <= 8'h00;
                15'h7664: d <= 8'h00; 15'h7665: d <= 8'h00; 15'h7666: d <= 8'h00; 15'h7667: d <= 8'h00;
                15'h7668: d <= 8'h00; 15'h7669: d <= 8'h00; 15'h766A: d <= 8'h00; 15'h766B: d <= 8'h00;
                15'h766C: d <= 8'h00; 15'h766D: d <= 8'h00; 15'h766E: d <= 8'h00; 15'h766F: d <= 8'h00;
                15'h7670: d <= 8'h00; 15'h7671: d <= 8'h00; 15'h7672: d <= 8'h00; 15'h7673: d <= 8'h00;
                15'h7674: d <= 8'h00; 15'h7675: d <= 8'h00; 15'h7676: d <= 8'h00; 15'h7677: d <= 8'h00;
                15'h7678: d <= 8'h00; 15'h7679: d <= 8'h00; 15'h767A: d <= 8'h00; 15'h767B: d <= 8'h00;
                15'h767C: d <= 8'h00; 15'h767D: d <= 8'h00; 15'h767E: d <= 8'h00; 15'h767F: d <= 8'hE0;
                15'h7680: d <= 8'h10; 15'h7681: d <= 8'h15; 15'h7682: d <= 8'h1A; 15'h7683: d <= 8'h1F;
                15'h7684: d <= 8'h20; 15'h7685: d <= 8'h25; 15'h7686: d <= 8'h2A; 15'h7687: d <= 8'h2F;
                15'h7688: d <= 8'h34; 15'h7689: d <= 8'h38; 15'h768A: d <= 8'h3C; 15'h768B: d <= 8'h31;
                15'h768C: d <= 8'h39; 15'h768D: d <= 8'h3D; 15'h768E: d <= 8'h32; 15'h768F: d <= 8'h36;
                15'h7690: d <= 8'h3E; 15'h7691: d <= 8'h33; 15'h7692: d <= 8'h37; 15'h7693: d <= 8'h3B;
                15'h7694: d <= 8'h44; 15'h7695: d <= 8'h48; 15'h7696: d <= 8'h4C; 15'h7697: d <= 8'h41;
                15'h7698: d <= 8'h49; 15'h7699: d <= 8'h4D; 15'h769A: d <= 8'h42; 15'h769B: d <= 8'h46;
                15'h769C: d <= 8'h4E; 15'h769D: d <= 8'h43; 15'h769E: d <= 8'h47; 15'h769F: d <= 8'h4B;
                15'h76A0: d <= 8'h50; 15'h76A1: d <= 8'h55; 15'h76A2: d <= 8'h5A; 15'h76A3: d <= 8'h5F;
                15'h76A4: d <= 8'h60; 15'h76A5: d <= 8'h65; 15'h76A6: d <= 8'h6A; 15'h76A7: d <= 8'h6F;
                15'h76A8: d <= 8'h74; 15'h76A9: d <= 8'h78; 15'h76AA: d <= 8'h7C; 15'h76AB: d <= 8'h71;
                15'h76AC: d <= 8'h79; 15'h76AD: d <= 8'h7D; 15'h76AE: d <= 8'h72; 15'h76AF: d <= 8'h76;
                15'h76B0: d <= 8'h7E; 15'h76B1: d <= 8'h73; 15'h76B2: d <= 8'h77; 15'h76B3: d <= 8'h7B;
                15'h76B4: d <= 8'h84; 15'h76B5: d <= 8'h88; 15'h76B6: d <= 8'h8C; 15'h76B7: d <= 8'h81;
                15'h76B8: d <= 8'h89; 15'h76B9: d <= 8'h8D; 15'h76BA: d <= 8'h82; 15'h76BB: d <= 8'h86;
                15'h76BC: d <= 8'h8E; 15'h76BD: d <= 8'h83; 15'h76BE: d <= 8'h87; 15'h76BF: d <= 8'h8B;
                15'h76C0: d <= 8'h90; 15'h76C1: d <= 8'h95; 15'h76C2: d <= 8'h9A; 15'h76C3: d <= 8'h9F;
                15'h76C4: d <= 8'hA4; 15'h76C5: d <= 8'hA8; 15'h76C6: d <= 8'hAC; 15'h76C7: d <= 8'hA1;
                15'h76C8: d <= 8'hA9; 15'h76C9: d <= 8'hAD; 15'h76CA: d <= 8'hA2; 15'h76CB: d <= 8'hA6;
                15'h76CC: d <= 8'hAE; 15'h76CD: d <= 8'hA3; 15'h76CE: d <= 8'hA7; 15'h76CF: d <= 8'hAB;
                15'h76D0: d <= 8'hB4; 15'h76D1: d <= 8'hB8; 15'h76D2: d <= 8'hBC; 15'h76D3: d <= 8'hB1;
                15'h76D4: d <= 8'hB9; 15'h76D5: d <= 8'hBD; 15'h76D6: d <= 8'hB2; 15'h76D7: d <= 8'hB6;
                15'h76D8: d <= 8'hBE; 15'h76D9: d <= 8'hB3; 15'h76DA: d <= 8'hB7; 15'h76DB: d <= 8'hBB;
                15'h76DC: d <= 8'hC4; 15'h76DD: d <= 8'hC8; 15'h76DE: d <= 8'hCC; 15'h76DF: d <= 8'hC1;
                15'h76E0: d <= 8'hC9; 15'h76E1: d <= 8'hCD; 15'h76E2: d <= 8'hC2; 15'h76E3: d <= 8'hC6;
                15'h76E4: d <= 8'hCE; 15'h76E5: d <= 8'hC3; 15'h76E6: d <= 8'hC7; 15'h76E7: d <= 8'hCB;
                15'h76E8: d <= 8'hC0; 15'h76E9: d <= 8'hC5; 15'h76EA: d <= 8'hCA; 15'h76EB: d <= 8'hCF;
                15'h76EC: d <= 8'hD0; 15'h76ED: d <= 8'hD5; 15'h76EE: d <= 8'hDA; 15'h76EF: d <= 8'hDF;
                15'h76F0: d <= 8'h74; 15'h76F1: d <= 8'h78; 15'h76F2: d <= 8'h7C; 15'h76F3: d <= 8'h71;
                15'h76F4: d <= 8'h79; 15'h76F5: d <= 8'h7D; 15'h76F6: d <= 8'h72; 15'h76F7: d <= 8'h76;
                15'h76F8: d <= 8'h7E; 15'h76F9: d <= 8'h73; 15'h76FA: d <= 8'h77; 15'h76FB: d <= 8'h7B;
                15'h76FC: d <= 8'hA0; 15'h76FD: d <= 8'hA5; 15'h76FE: d <= 8'hAA; 15'h76FF: d <= 8'hAF;
                15'h7700: d <= 8'h00; 15'h7701: d <= 8'h00; 15'h7702: d <= 8'h00; 15'h7703: d <= 8'h00;
                15'h7704: d <= 8'h00; 15'h7705: d <= 8'h00; 15'h7706: d <= 8'h00; 15'h7707: d <= 8'h00;
                15'h7708: d <= 8'h00; 15'h7709: d <= 8'h00; 15'h770A: d <= 8'h00; 15'h770B: d <= 8'h00;
                15'h770C: d <= 8'h00; 15'h770D: d <= 8'h00; 15'h770E: d <= 8'h00; 15'h770F: d <= 8'h00;
                15'h7710: d <= 8'h00; 15'h7711: d <= 8'h00; 15'h7712: d <= 8'h00; 15'h7713: d <= 8'h00;
                15'h7714: d <= 8'h00; 15'h7715: d <= 8'h00; 15'h7716: d <= 8'h00; 15'h7717: d <= 8'h00;
                15'h7718: d <= 8'h00; 15'h7719: d <= 8'h00; 15'h771A: d <= 8'h00; 15'h771B: d <= 8'h00;
                15'h771C: d <= 8'h00; 15'h771D: d <= 8'h00; 15'h771E: d <= 8'h00; 15'h771F: d <= 8'h00;
                15'h7720: d <= 8'h00; 15'h7721: d <= 8'h00; 15'h7722: d <= 8'h00; 15'h7723: d <= 8'h00;
                15'h7724: d <= 8'h00; 15'h7725: d <= 8'h00; 15'h7726: d <= 8'h00; 15'h7727: d <= 8'h00;
                15'h7728: d <= 8'h00; 15'h7729: d <= 8'h00; 15'h772A: d <= 8'h00; 15'h772B: d <= 8'h00;
                15'h772C: d <= 8'h00; 15'h772D: d <= 8'h00; 15'h772E: d <= 8'h00; 15'h772F: d <= 8'hAF;
                15'h7730: d <= 8'h00; 15'h7731: d <= 8'h00; 15'h7732: d <= 8'h00; 15'h7733: d <= 8'h00;
                15'h7734: d <= 8'h00; 15'h7735: d <= 8'h00; 15'h7736: d <= 8'h00; 15'h7737: d <= 8'h00;
                15'h7738: d <= 8'h00; 15'h7739: d <= 8'h00; 15'h773A: d <= 8'h00; 15'h773B: d <= 8'h00;
                15'h773C: d <= 8'h00; 15'h773D: d <= 8'h00; 15'h773E: d <= 8'h00; 15'h773F: d <= 8'h00;
                15'h7740: d <= 8'h00; 15'h7741: d <= 8'h00; 15'h7742: d <= 8'h00; 15'h7743: d <= 8'h00;
                15'h7744: d <= 8'h00; 15'h7745: d <= 8'h00; 15'h7746: d <= 8'h00; 15'h7747: d <= 8'h00;
                15'h7748: d <= 8'h00; 15'h7749: d <= 8'h00; 15'h774A: d <= 8'h00; 15'h774B: d <= 8'h00;
                15'h774C: d <= 8'h00; 15'h774D: d <= 8'h00; 15'h774E: d <= 8'h00; 15'h774F: d <= 8'h00;
                15'h7750: d <= 8'h00; 15'h7751: d <= 8'h00; 15'h7752: d <= 8'h00; 15'h7753: d <= 8'h00;
                15'h7754: d <= 8'h00; 15'h7755: d <= 8'h00; 15'h7756: d <= 8'h00; 15'h7757: d <= 8'h00;
                15'h7758: d <= 8'h45; 15'h7759: d <= 8'h35; 15'h775A: d <= 8'hAA; 15'h775B: d <= 8'h00;
                15'h775C: d <= 8'h00; 15'h775D: d <= 8'h00; 15'h775E: d <= 8'h00; 15'h775F: d <= 8'h00;
                15'h7760: d <= 8'h00; 15'h7761: d <= 8'h00; 15'h7762: d <= 8'h00; 15'h7763: d <= 8'h00;
                15'h7764: d <= 8'h00; 15'h7765: d <= 8'h00; 15'h7766: d <= 8'h00; 15'h7767: d <= 8'h00;
                15'h7768: d <= 8'h00; 15'h7769: d <= 8'h00; 15'h776A: d <= 8'h00; 15'h776B: d <= 8'h00;
                15'h776C: d <= 8'h00; 15'h776D: d <= 8'h00; 15'h776E: d <= 8'h00; 15'h776F: d <= 8'h00;
                15'h7770: d <= 8'h00; 15'h7771: d <= 8'h00; 15'h7772: d <= 8'h00; 15'h7773: d <= 8'h00;
                15'h7774: d <= 8'h00; 15'h7775: d <= 8'h00; 15'h7776: d <= 8'h00; 15'h7777: d <= 8'h00;
                15'h7778: d <= 8'h00; 15'h7779: d <= 8'h00; 15'h777A: d <= 8'h00; 15'h777B: d <= 8'h00;
                15'h777C: d <= 8'h00; 15'h777D: d <= 8'h00; 15'h777E: d <= 8'h00; 15'h777F: d <= 8'hE0;
                15'h7780: d <= 8'h10; 15'h7781: d <= 8'h15; 15'h7782: d <= 8'h1A; 15'h7783: d <= 8'h1F;
                15'h7784: d <= 8'h20; 15'h7785: d <= 8'h25; 15'h7786: d <= 8'h2A; 15'h7787: d <= 8'h2F;
                15'h7788: d <= 8'h34; 15'h7789: d <= 8'h38; 15'h778A: d <= 8'h3C; 15'h778B: d <= 8'h31;
                15'h778C: d <= 8'h39; 15'h778D: d <= 8'h3D; 15'h778E: d <= 8'h32; 15'h778F: d <= 8'h36;
                15'h7790: d <= 8'h3E; 15'h7791: d <= 8'h33; 15'h7792: d <= 8'h37; 15'h7793: d <= 8'h3B;
                15'h7794: d <= 8'h44; 15'h7795: d <= 8'h48; 15'h7796: d <= 8'h4C; 15'h7797: d <= 8'h41;
                15'h7798: d <= 8'h49; 15'h7799: d <= 8'h4D; 15'h779A: d <= 8'h42; 15'h779B: d <= 8'h46;
                15'h779C: d <= 8'h4E; 15'h779D: d <= 8'h43; 15'h779E: d <= 8'h47; 15'h779F: d <= 8'h4B;
                15'h77A0: d <= 8'h50; 15'h77A1: d <= 8'h55; 15'h77A2: d <= 8'h5A; 15'h77A3: d <= 8'h5F;
                15'h77A4: d <= 8'h60; 15'h77A5: d <= 8'h65; 15'h77A6: d <= 8'h6A; 15'h77A7: d <= 8'h6F;
                15'h77A8: d <= 8'h74; 15'h77A9: d <= 8'h78; 15'h77AA: d <= 8'h7C; 15'h77AB: d <= 8'h71;
                15'h77AC: d <= 8'h79; 15'h77AD: d <= 8'h7D; 15'h77AE: d <= 8'h72; 15'h77AF: d <= 8'h76;
                15'h77B0: d <= 8'h7E; 15'h77B1: d <= 8'h73; 15'h77B2: d <= 8'h77; 15'h77B3: d <= 8'h7B;
                15'h77B4: d <= 8'h84; 15'h77B5: d <= 8'h88; 15'h77B6: d <= 8'h8C; 15'h77B7: d <= 8'h81;
                15'h77B8: d <= 8'h89; 15'h77B9: d <= 8'h8D; 15'h77BA: d <= 8'h82; 15'h77BB: d <= 8'h86;
                15'h77BC: d <= 8'h8E; 15'h77BD: d <= 8'h83; 15'h77BE: d <= 8'h87; 15'h77BF: d <= 8'h8B;
                15'h77C0: d <= 8'h90; 15'h77C1: d <= 8'h95; 15'h77C2: d <= 8'h9A; 15'h77C3: d <= 8'h9F;
                15'h77C4: d <= 8'hA4; 15'h77C5: d <= 8'hA8; 15'h77C6: d <= 8'hAC; 15'h77C7: d <= 8'hA1;
                15'h77C8: d <= 8'hA9; 15'h77C9: d <= 8'hAD; 15'h77CA: d <= 8'hA2; 15'h77CB: d <= 8'hA6;
                15'h77CC: d <= 8'hAE; 15'h77CD: d <= 8'hA3; 15'h77CE: d <= 8'hA7; 15'h77CF: d <= 8'hAB;
                15'h77D0: d <= 8'hB4; 15'h77D1: d <= 8'hB8; 15'h77D2: d <= 8'hBC; 15'h77D3: d <= 8'hB1;
                15'h77D4: d <= 8'hB9; 15'h77D5: d <= 8'hBD; 15'h77D6: d <= 8'hB2; 15'h77D7: d <= 8'hB6;
                15'h77D8: d <= 8'hBE; 15'h77D9: d <= 8'hB3; 15'h77DA: d <= 8'hB7; 15'h77DB: d <= 8'hBB;
                15'h77DC: d <= 8'hC4; 15'h77DD: d <= 8'hC8; 15'h77DE: d <= 8'hCC; 15'h77DF: d <= 8'hC1;
                15'h77E0: d <= 8'hC9; 15'h77E1: d <= 8'hCD; 15'h77E2: d <= 8'hC2; 15'h77E3: d <= 8'hC6;
                15'h77E4: d <= 8'hCE; 15'h77E5: d <= 8'hC3; 15'h77E6: d <= 8'hC7; 15'h77E7: d <= 8'hCB;
                15'h77E8: d <= 8'hC0; 15'h77E9: d <= 8'hC5; 15'h77EA: d <= 8'hCA; 15'h77EB: d <= 8'hCF;
                15'h77EC: d <= 8'hD0; 15'h77ED: d <= 8'hD5; 15'h77EE: d <= 8'hDA; 15'h77EF: d <= 8'hDF;
                15'h77F0: d <= 8'h74; 15'h77F1: d <= 8'h78; 15'h77F2: d <= 8'h7C; 15'h77F3: d <= 8'h71;
                15'h77F4: d <= 8'h79; 15'h77F5: d <= 8'h7D; 15'h77F6: d <= 8'h72; 15'h77F7: d <= 8'h76;
                15'h77F8: d <= 8'h7E; 15'h77F9: d <= 8'h73; 15'h77FA: d <= 8'h77; 15'h77FB: d <= 8'h7B;
                15'h77FC: d <= 8'hA0; 15'h77FD: d <= 8'hA5; 15'h77FE: d <= 8'hAA; 15'h77FF: d <= 8'hAF;
                15'h7800: d <= 8'h00; 15'h7801: d <= 8'h00; 15'h7802: d <= 8'h00; 15'h7803: d <= 8'h00;
                15'h7804: d <= 8'h00; 15'h7805: d <= 8'h00; 15'h7806: d <= 8'h00; 15'h7807: d <= 8'h00;
                15'h7808: d <= 8'h00; 15'h7809: d <= 8'h00; 15'h780A: d <= 8'h00; 15'h780B: d <= 8'h00;
                15'h780C: d <= 8'h00; 15'h780D: d <= 8'h00; 15'h780E: d <= 8'h00; 15'h780F: d <= 8'h00;
                15'h7810: d <= 8'h00; 15'h7811: d <= 8'h00; 15'h7812: d <= 8'h00; 15'h7813: d <= 8'h00;
                15'h7814: d <= 8'h00; 15'h7815: d <= 8'h00; 15'h7816: d <= 8'h00; 15'h7817: d <= 8'h00;
                15'h7818: d <= 8'h00; 15'h7819: d <= 8'h00; 15'h781A: d <= 8'h00; 15'h781B: d <= 8'h00;
                15'h781C: d <= 8'h00; 15'h781D: d <= 8'h00; 15'h781E: d <= 8'h00; 15'h781F: d <= 8'h00;
                15'h7820: d <= 8'h00; 15'h7821: d <= 8'h00; 15'h7822: d <= 8'h00; 15'h7823: d <= 8'h00;
                15'h7824: d <= 8'h00; 15'h7825: d <= 8'h00; 15'h7826: d <= 8'h00; 15'h7827: d <= 8'h00;
                15'h7828: d <= 8'h00; 15'h7829: d <= 8'h00; 15'h782A: d <= 8'h00; 15'h782B: d <= 8'h00;
                15'h782C: d <= 8'h00; 15'h782D: d <= 8'h00; 15'h782E: d <= 8'h00; 15'h782F: d <= 8'h7B;
                15'h7830: d <= 8'h00; 15'h7831: d <= 8'h00; 15'h7832: d <= 8'h00; 15'h7833: d <= 8'h00;
                15'h7834: d <= 8'h00; 15'h7835: d <= 8'h00; 15'h7836: d <= 8'h00; 15'h7837: d <= 8'h00;
                15'h7838: d <= 8'h00; 15'h7839: d <= 8'h00; 15'h783A: d <= 8'h00; 15'h783B: d <= 8'h00;
                15'h783C: d <= 8'h00; 15'h783D: d <= 8'h00; 15'h783E: d <= 8'h00; 15'h783F: d <= 8'h00;
                15'h7840: d <= 8'h00; 15'h7841: d <= 8'h00; 15'h7842: d <= 8'h00; 15'h7843: d <= 8'h00;
                15'h7844: d <= 8'h00; 15'h7845: d <= 8'h00; 15'h7846: d <= 8'h00; 15'h7847: d <= 8'h00;
                15'h7848: d <= 8'h00; 15'h7849: d <= 8'h00; 15'h784A: d <= 8'h00; 15'h784B: d <= 8'h00;
                15'h784C: d <= 8'h00; 15'h784D: d <= 8'h00; 15'h784E: d <= 8'h00; 15'h784F: d <= 8'h00;
                15'h7850: d <= 8'h00; 15'h7851: d <= 8'h00; 15'h7852: d <= 8'h00; 15'h7853: d <= 8'h00;
                15'h7854: d <= 8'h00; 15'h7855: d <= 8'h00; 15'h7856: d <= 8'h00; 15'h7857: d <= 8'h00;
                15'h7858: d <= 8'h45; 15'h7859: d <= 8'h35; 15'h785A: d <= 8'h32; 15'h785B: d <= 8'h00;
                15'h785C: d <= 8'h00; 15'h785D: d <= 8'h00; 15'h785E: d <= 8'h00; 15'h785F: d <= 8'h00;
                15'h7860: d <= 8'h00; 15'h7861: d <= 8'h00; 15'h7862: d <= 8'h00; 15'h7863: d <= 8'h00;
                15'h7864: d <= 8'h00; 15'h7865: d <= 8'h00; 15'h7866: d <= 8'h00; 15'h7867: d <= 8'h00;
                15'h7868: d <= 8'h00; 15'h7869: d <= 8'h00; 15'h786A: d <= 8'h00; 15'h786B: d <= 8'h00;
                15'h786C: d <= 8'h00; 15'h786D: d <= 8'h00; 15'h786E: d <= 8'h00; 15'h786F: d <= 8'h00;
                15'h7870: d <= 8'h00; 15'h7871: d <= 8'h00; 15'h7872: d <= 8'h00; 15'h7873: d <= 8'h00;
                15'h7874: d <= 8'h00; 15'h7875: d <= 8'h00; 15'h7876: d <= 8'h00; 15'h7877: d <= 8'h00;
                15'h7878: d <= 8'h00; 15'h7879: d <= 8'h00; 15'h787A: d <= 8'h00; 15'h787B: d <= 8'h00;
                15'h787C: d <= 8'h00; 15'h787D: d <= 8'h00; 15'h787E: d <= 8'h00; 15'h787F: d <= 8'hE0;
                15'h7880: d <= 8'h10; 15'h7881: d <= 8'h15; 15'h7882: d <= 8'h1A; 15'h7883: d <= 8'h1F;
                15'h7884: d <= 8'h20; 15'h7885: d <= 8'h25; 15'h7886: d <= 8'h2A; 15'h7887: d <= 8'h2F;
                15'h7888: d <= 8'h34; 15'h7889: d <= 8'h38; 15'h788A: d <= 8'h3C; 15'h788B: d <= 8'h31;
                15'h788C: d <= 8'h39; 15'h788D: d <= 8'h3D; 15'h788E: d <= 8'h32; 15'h788F: d <= 8'h36;
                15'h7890: d <= 8'h3E; 15'h7891: d <= 8'h33; 15'h7892: d <= 8'h37; 15'h7893: d <= 8'h3B;
                15'h7894: d <= 8'h44; 15'h7895: d <= 8'h48; 15'h7896: d <= 8'h4C; 15'h7897: d <= 8'h41;
                15'h7898: d <= 8'h49; 15'h7899: d <= 8'h4D; 15'h789A: d <= 8'h42; 15'h789B: d <= 8'h46;
                15'h789C: d <= 8'h4E; 15'h789D: d <= 8'h43; 15'h789E: d <= 8'h47; 15'h789F: d <= 8'h4B;
                15'h78A0: d <= 8'h50; 15'h78A1: d <= 8'h55; 15'h78A2: d <= 8'h5A; 15'h78A3: d <= 8'h5F;
                15'h78A4: d <= 8'h60; 15'h78A5: d <= 8'h65; 15'h78A6: d <= 8'h6A; 15'h78A7: d <= 8'h6F;
                15'h78A8: d <= 8'h74; 15'h78A9: d <= 8'h78; 15'h78AA: d <= 8'h7C; 15'h78AB: d <= 8'h71;
                15'h78AC: d <= 8'h79; 15'h78AD: d <= 8'h7D; 15'h78AE: d <= 8'h72; 15'h78AF: d <= 8'h76;
                15'h78B0: d <= 8'h7E; 15'h78B1: d <= 8'h73; 15'h78B2: d <= 8'h77; 15'h78B3: d <= 8'h7B;
                15'h78B4: d <= 8'h84; 15'h78B5: d <= 8'h88; 15'h78B6: d <= 8'h8C; 15'h78B7: d <= 8'h81;
                15'h78B8: d <= 8'h89; 15'h78B9: d <= 8'h8D; 15'h78BA: d <= 8'h82; 15'h78BB: d <= 8'h86;
                15'h78BC: d <= 8'h8E; 15'h78BD: d <= 8'h83; 15'h78BE: d <= 8'h87; 15'h78BF: d <= 8'h8B;
                15'h78C0: d <= 8'h90; 15'h78C1: d <= 8'h95; 15'h78C2: d <= 8'h9A; 15'h78C3: d <= 8'h9F;
                15'h78C4: d <= 8'hA4; 15'h78C5: d <= 8'hA8; 15'h78C6: d <= 8'hAC; 15'h78C7: d <= 8'hA1;
                15'h78C8: d <= 8'hA9; 15'h78C9: d <= 8'hAD; 15'h78CA: d <= 8'hA2; 15'h78CB: d <= 8'hA6;
                15'h78CC: d <= 8'hAE; 15'h78CD: d <= 8'hA3; 15'h78CE: d <= 8'hA7; 15'h78CF: d <= 8'hAB;
                15'h78D0: d <= 8'hB4; 15'h78D1: d <= 8'hB8; 15'h78D2: d <= 8'hBC; 15'h78D3: d <= 8'hB1;
                15'h78D4: d <= 8'hB9; 15'h78D5: d <= 8'hBD; 15'h78D6: d <= 8'hB2; 15'h78D7: d <= 8'hB6;
                15'h78D8: d <= 8'hBE; 15'h78D9: d <= 8'hB3; 15'h78DA: d <= 8'hB7; 15'h78DB: d <= 8'hBB;
                15'h78DC: d <= 8'hC4; 15'h78DD: d <= 8'hC8; 15'h78DE: d <= 8'hCC; 15'h78DF: d <= 8'hC1;
                15'h78E0: d <= 8'hC9; 15'h78E1: d <= 8'hCD; 15'h78E2: d <= 8'hC2; 15'h78E3: d <= 8'hC6;
                15'h78E4: d <= 8'hCE; 15'h78E5: d <= 8'hC3; 15'h78E6: d <= 8'hC7; 15'h78E7: d <= 8'hCB;
                15'h78E8: d <= 8'hC0; 15'h78E9: d <= 8'hC5; 15'h78EA: d <= 8'hCA; 15'h78EB: d <= 8'hCF;
                15'h78EC: d <= 8'hD0; 15'h78ED: d <= 8'hD5; 15'h78EE: d <= 8'hDA; 15'h78EF: d <= 8'hDF;
                15'h78F0: d <= 8'h74; 15'h78F1: d <= 8'h78; 15'h78F2: d <= 8'h7C; 15'h78F3: d <= 8'h71;
                15'h78F4: d <= 8'h79; 15'h78F5: d <= 8'h7D; 15'h78F6: d <= 8'h72; 15'h78F7: d <= 8'h76;
                15'h78F8: d <= 8'h7E; 15'h78F9: d <= 8'h73; 15'h78FA: d <= 8'h77; 15'h78FB: d <= 8'h7B;
                15'h78FC: d <= 8'hA0; 15'h78FD: d <= 8'hA5; 15'h78FE: d <= 8'hAA; 15'h78FF: d <= 8'hAF;
                15'h7900: d <= 8'h00; 15'h7901: d <= 8'h00; 15'h7902: d <= 8'h00; 15'h7903: d <= 8'h00;
                15'h7904: d <= 8'h00; 15'h7905: d <= 8'h00; 15'h7906: d <= 8'h00; 15'h7907: d <= 8'h00;
                15'h7908: d <= 8'h00; 15'h7909: d <= 8'h00; 15'h790A: d <= 8'h00; 15'h790B: d <= 8'h00;
                15'h790C: d <= 8'h00; 15'h790D: d <= 8'h00; 15'h790E: d <= 8'h00; 15'h790F: d <= 8'h00;
                15'h7910: d <= 8'h00; 15'h7911: d <= 8'h00; 15'h7912: d <= 8'h00; 15'h7913: d <= 8'h00;
                15'h7914: d <= 8'h00; 15'h7915: d <= 8'h00; 15'h7916: d <= 8'h00; 15'h7917: d <= 8'h00;
                15'h7918: d <= 8'h00; 15'h7919: d <= 8'h00; 15'h791A: d <= 8'h00; 15'h791B: d <= 8'h00;
                15'h791C: d <= 8'h00; 15'h791D: d <= 8'h00; 15'h791E: d <= 8'h00; 15'h791F: d <= 8'h00;
                15'h7920: d <= 8'h00; 15'h7921: d <= 8'h00; 15'h7922: d <= 8'h00; 15'h7923: d <= 8'h00;
                15'h7924: d <= 8'h00; 15'h7925: d <= 8'h00; 15'h7926: d <= 8'h00; 15'h7927: d <= 8'h00;
                15'h7928: d <= 8'h00; 15'h7929: d <= 8'h00; 15'h792A: d <= 8'h00; 15'h792B: d <= 8'h00;
                15'h792C: d <= 8'h00; 15'h792D: d <= 8'h00; 15'h792E: d <= 8'h00; 15'h792F: d <= 8'h7B;
                15'h7930: d <= 8'h00; 15'h7931: d <= 8'h00; 15'h7932: d <= 8'h00; 15'h7933: d <= 8'h00;
                15'h7934: d <= 8'h00; 15'h7935: d <= 8'h00; 15'h7936: d <= 8'h00; 15'h7937: d <= 8'h00;
                15'h7938: d <= 8'h00; 15'h7939: d <= 8'h00; 15'h793A: d <= 8'h00; 15'h793B: d <= 8'h00;
                15'h793C: d <= 8'h00; 15'h793D: d <= 8'h00; 15'h793E: d <= 8'h00; 15'h793F: d <= 8'h00;
                15'h7940: d <= 8'h00; 15'h7941: d <= 8'h00; 15'h7942: d <= 8'h00; 15'h7943: d <= 8'h00;
                15'h7944: d <= 8'h00; 15'h7945: d <= 8'h00; 15'h7946: d <= 8'h00; 15'h7947: d <= 8'h00;
                15'h7948: d <= 8'h00; 15'h7949: d <= 8'h00; 15'h794A: d <= 8'h00; 15'h794B: d <= 8'h00;
                15'h794C: d <= 8'h00; 15'h794D: d <= 8'h00; 15'h794E: d <= 8'h00; 15'h794F: d <= 8'h00;
                15'h7950: d <= 8'h00; 15'h7951: d <= 8'h00; 15'h7952: d <= 8'h00; 15'h7953: d <= 8'h00;
                15'h7954: d <= 8'h00; 15'h7955: d <= 8'h00; 15'h7956: d <= 8'h00; 15'h7957: d <= 8'h00;
                15'h7958: d <= 8'h45; 15'h7959: d <= 8'h35; 15'h795A: d <= 8'h32; 15'h795B: d <= 8'h00;
                15'h795C: d <= 8'h00; 15'h795D: d <= 8'h00; 15'h795E: d <= 8'h00; 15'h795F: d <= 8'h00;
                15'h7960: d <= 8'h00; 15'h7961: d <= 8'h00; 15'h7962: d <= 8'h00; 15'h7963: d <= 8'h00;
                15'h7964: d <= 8'h00; 15'h7965: d <= 8'h00; 15'h7966: d <= 8'h00; 15'h7967: d <= 8'h00;
                15'h7968: d <= 8'h00; 15'h7969: d <= 8'h00; 15'h796A: d <= 8'h00; 15'h796B: d <= 8'h00;
                15'h796C: d <= 8'h00; 15'h796D: d <= 8'h00; 15'h796E: d <= 8'h00; 15'h796F: d <= 8'h00;
                15'h7970: d <= 8'h00; 15'h7971: d <= 8'h00; 15'h7972: d <= 8'h00; 15'h7973: d <= 8'h00;
                15'h7974: d <= 8'h00; 15'h7975: d <= 8'h00; 15'h7976: d <= 8'h00; 15'h7977: d <= 8'h00;
                15'h7978: d <= 8'h00; 15'h7979: d <= 8'h00; 15'h797A: d <= 8'h00; 15'h797B: d <= 8'h00;
                15'h797C: d <= 8'h00; 15'h797D: d <= 8'h00; 15'h797E: d <= 8'h00; 15'h797F: d <= 8'hE0;
                15'h7980: d <= 8'h10; 15'h7981: d <= 8'h15; 15'h7982: d <= 8'h1A; 15'h7983: d <= 8'h1F;
                15'h7984: d <= 8'h20; 15'h7985: d <= 8'h25; 15'h7986: d <= 8'h2A; 15'h7987: d <= 8'h2F;
                15'h7988: d <= 8'h34; 15'h7989: d <= 8'h38; 15'h798A: d <= 8'h3C; 15'h798B: d <= 8'h31;
                15'h798C: d <= 8'h39; 15'h798D: d <= 8'h3D; 15'h798E: d <= 8'h32; 15'h798F: d <= 8'h36;
                15'h7990: d <= 8'h3E; 15'h7991: d <= 8'h33; 15'h7992: d <= 8'h37; 15'h7993: d <= 8'h3B;
                15'h7994: d <= 8'h44; 15'h7995: d <= 8'h48; 15'h7996: d <= 8'h4C; 15'h7997: d <= 8'h41;
                15'h7998: d <= 8'h49; 15'h7999: d <= 8'h4D; 15'h799A: d <= 8'h42; 15'h799B: d <= 8'h46;
                15'h799C: d <= 8'h4E; 15'h799D: d <= 8'h43; 15'h799E: d <= 8'h47; 15'h799F: d <= 8'h4B;
                15'h79A0: d <= 8'h50; 15'h79A1: d <= 8'h55; 15'h79A2: d <= 8'h5A; 15'h79A3: d <= 8'h5F;
                15'h79A4: d <= 8'h60; 15'h79A5: d <= 8'h65; 15'h79A6: d <= 8'h6A; 15'h79A7: d <= 8'h6F;
                15'h79A8: d <= 8'h74; 15'h79A9: d <= 8'h78; 15'h79AA: d <= 8'h7C; 15'h79AB: d <= 8'h71;
                15'h79AC: d <= 8'h79; 15'h79AD: d <= 8'h7D; 15'h79AE: d <= 8'h72; 15'h79AF: d <= 8'h76;
                15'h79B0: d <= 8'h7E; 15'h79B1: d <= 8'h73; 15'h79B2: d <= 8'h77; 15'h79B3: d <= 8'h7B;
                15'h79B4: d <= 8'h84; 15'h79B5: d <= 8'h88; 15'h79B6: d <= 8'h8C; 15'h79B7: d <= 8'h81;
                15'h79B8: d <= 8'h89; 15'h79B9: d <= 8'h8D; 15'h79BA: d <= 8'h82; 15'h79BB: d <= 8'h86;
                15'h79BC: d <= 8'h8E; 15'h79BD: d <= 8'h83; 15'h79BE: d <= 8'h87; 15'h79BF: d <= 8'h8B;
                15'h79C0: d <= 8'h90; 15'h79C1: d <= 8'h95; 15'h79C2: d <= 8'h9A; 15'h79C3: d <= 8'h9F;
                15'h79C4: d <= 8'hA4; 15'h79C5: d <= 8'hA8; 15'h79C6: d <= 8'hAC; 15'h79C7: d <= 8'hA1;
                15'h79C8: d <= 8'hA9; 15'h79C9: d <= 8'hAD; 15'h79CA: d <= 8'hA2; 15'h79CB: d <= 8'hA6;
                15'h79CC: d <= 8'hAE; 15'h79CD: d <= 8'hA3; 15'h79CE: d <= 8'hA7; 15'h79CF: d <= 8'hAB;
                15'h79D0: d <= 8'hB4; 15'h79D1: d <= 8'hB8; 15'h79D2: d <= 8'hBC; 15'h79D3: d <= 8'hB1;
                15'h79D4: d <= 8'hB9; 15'h79D5: d <= 8'hBD; 15'h79D6: d <= 8'hB2; 15'h79D7: d <= 8'hB6;
                15'h79D8: d <= 8'hBE; 15'h79D9: d <= 8'hB3; 15'h79DA: d <= 8'hB7; 15'h79DB: d <= 8'hBB;
                15'h79DC: d <= 8'hC4; 15'h79DD: d <= 8'hC8; 15'h79DE: d <= 8'hCC; 15'h79DF: d <= 8'hC1;
                15'h79E0: d <= 8'hC9; 15'h79E1: d <= 8'hCD; 15'h79E2: d <= 8'hC2; 15'h79E3: d <= 8'hC6;
                15'h79E4: d <= 8'hCE; 15'h79E5: d <= 8'hC3; 15'h79E6: d <= 8'hC7; 15'h79E7: d <= 8'hCB;
                15'h79E8: d <= 8'hC0; 15'h79E9: d <= 8'hC5; 15'h79EA: d <= 8'hCA; 15'h79EB: d <= 8'hCF;
                15'h79EC: d <= 8'hD0; 15'h79ED: d <= 8'hD5; 15'h79EE: d <= 8'hDA; 15'h79EF: d <= 8'hDF;
                15'h79F0: d <= 8'h74; 15'h79F1: d <= 8'h78; 15'h79F2: d <= 8'h7C; 15'h79F3: d <= 8'h71;
                15'h79F4: d <= 8'h79; 15'h79F5: d <= 8'h7D; 15'h79F6: d <= 8'h72; 15'h79F7: d <= 8'h76;
                15'h79F8: d <= 8'h7E; 15'h79F9: d <= 8'h73; 15'h79FA: d <= 8'h77; 15'h79FB: d <= 8'h7B;
                15'h79FC: d <= 8'hA0; 15'h79FD: d <= 8'hA5; 15'h79FE: d <= 8'hAA; 15'h79FF: d <= 8'hAF;
                15'h7A00: d <= 8'h00; 15'h7A01: d <= 8'h00; 15'h7A02: d <= 8'h00; 15'h7A03: d <= 8'h00;
                15'h7A04: d <= 8'h00; 15'h7A05: d <= 8'h00; 15'h7A06: d <= 8'h00; 15'h7A07: d <= 8'h00;
                15'h7A08: d <= 8'h00; 15'h7A09: d <= 8'h00; 15'h7A0A: d <= 8'h00; 15'h7A0B: d <= 8'h00;
                15'h7A0C: d <= 8'h00; 15'h7A0D: d <= 8'h00; 15'h7A0E: d <= 8'h00; 15'h7A0F: d <= 8'h00;
                15'h7A10: d <= 8'h00; 15'h7A11: d <= 8'h00; 15'h7A12: d <= 8'h00; 15'h7A13: d <= 8'h00;
                15'h7A14: d <= 8'h00; 15'h7A15: d <= 8'h00; 15'h7A16: d <= 8'h00; 15'h7A17: d <= 8'h00;
                15'h7A18: d <= 8'h00; 15'h7A19: d <= 8'h00; 15'h7A1A: d <= 8'h00; 15'h7A1B: d <= 8'h00;
                15'h7A1C: d <= 8'h00; 15'h7A1D: d <= 8'h00; 15'h7A1E: d <= 8'h00; 15'h7A1F: d <= 8'h00;
                15'h7A20: d <= 8'h00; 15'h7A21: d <= 8'h00; 15'h7A22: d <= 8'h00; 15'h7A23: d <= 8'h00;
                15'h7A24: d <= 8'h00; 15'h7A25: d <= 8'h00; 15'h7A26: d <= 8'h00; 15'h7A27: d <= 8'h00;
                15'h7A28: d <= 8'h00; 15'h7A29: d <= 8'h00; 15'h7A2A: d <= 8'h00; 15'h7A2B: d <= 8'h00;
                15'h7A2C: d <= 8'h00; 15'h7A2D: d <= 8'h00; 15'h7A2E: d <= 8'h00; 15'h7A2F: d <= 8'h7B;
                15'h7A30: d <= 8'h00; 15'h7A31: d <= 8'h00; 15'h7A32: d <= 8'h00; 15'h7A33: d <= 8'h00;
                15'h7A34: d <= 8'h00; 15'h7A35: d <= 8'h00; 15'h7A36: d <= 8'h00; 15'h7A37: d <= 8'h00;
                15'h7A38: d <= 8'h00; 15'h7A39: d <= 8'h00; 15'h7A3A: d <= 8'h00; 15'h7A3B: d <= 8'h00;
                15'h7A3C: d <= 8'h00; 15'h7A3D: d <= 8'h00; 15'h7A3E: d <= 8'h00; 15'h7A3F: d <= 8'h00;
                15'h7A40: d <= 8'h00; 15'h7A41: d <= 8'h00; 15'h7A42: d <= 8'h00; 15'h7A43: d <= 8'h00;
                15'h7A44: d <= 8'h00; 15'h7A45: d <= 8'h00; 15'h7A46: d <= 8'h00; 15'h7A47: d <= 8'h00;
                15'h7A48: d <= 8'h00; 15'h7A49: d <= 8'h00; 15'h7A4A: d <= 8'h00; 15'h7A4B: d <= 8'h00;
                15'h7A4C: d <= 8'h00; 15'h7A4D: d <= 8'h00; 15'h7A4E: d <= 8'h00; 15'h7A4F: d <= 8'h00;
                15'h7A50: d <= 8'h00; 15'h7A51: d <= 8'h00; 15'h7A52: d <= 8'h00; 15'h7A53: d <= 8'h00;
                15'h7A54: d <= 8'h00; 15'h7A55: d <= 8'h00; 15'h7A56: d <= 8'h00; 15'h7A57: d <= 8'h00;
                15'h7A58: d <= 8'h45; 15'h7A59: d <= 8'h35; 15'h7A5A: d <= 8'h32; 15'h7A5B: d <= 8'h00;
                15'h7A5C: d <= 8'h00; 15'h7A5D: d <= 8'h00; 15'h7A5E: d <= 8'h00; 15'h7A5F: d <= 8'h00;
                15'h7A60: d <= 8'h00; 15'h7A61: d <= 8'h00; 15'h7A62: d <= 8'h00; 15'h7A63: d <= 8'h00;
                15'h7A64: d <= 8'h00; 15'h7A65: d <= 8'h00; 15'h7A66: d <= 8'h00; 15'h7A67: d <= 8'h00;
                15'h7A68: d <= 8'h00; 15'h7A69: d <= 8'h00; 15'h7A6A: d <= 8'h00; 15'h7A6B: d <= 8'h00;
                15'h7A6C: d <= 8'h00; 15'h7A6D: d <= 8'h00; 15'h7A6E: d <= 8'h00; 15'h7A6F: d <= 8'h00;
                15'h7A70: d <= 8'h00; 15'h7A71: d <= 8'h00; 15'h7A72: d <= 8'h00; 15'h7A73: d <= 8'h00;
                15'h7A74: d <= 8'h00; 15'h7A75: d <= 8'h00; 15'h7A76: d <= 8'h00; 15'h7A77: d <= 8'h00;
                15'h7A78: d <= 8'h00; 15'h7A79: d <= 8'h00; 15'h7A7A: d <= 8'h00; 15'h7A7B: d <= 8'h00;
                15'h7A7C: d <= 8'h00; 15'h7A7D: d <= 8'h00; 15'h7A7E: d <= 8'h00; 15'h7A7F: d <= 8'hE0;
                15'h7A80: d <= 8'h10; 15'h7A81: d <= 8'h15; 15'h7A82: d <= 8'h1A; 15'h7A83: d <= 8'h1F;
                15'h7A84: d <= 8'h20; 15'h7A85: d <= 8'h25; 15'h7A86: d <= 8'h2A; 15'h7A87: d <= 8'h2F;
                15'h7A88: d <= 8'h34; 15'h7A89: d <= 8'h38; 15'h7A8A: d <= 8'h3C; 15'h7A8B: d <= 8'h31;
                15'h7A8C: d <= 8'h39; 15'h7A8D: d <= 8'h3D; 15'h7A8E: d <= 8'h32; 15'h7A8F: d <= 8'h36;
                15'h7A90: d <= 8'h3E; 15'h7A91: d <= 8'h33; 15'h7A92: d <= 8'h37; 15'h7A93: d <= 8'h3B;
                15'h7A94: d <= 8'h44; 15'h7A95: d <= 8'h48; 15'h7A96: d <= 8'h4C; 15'h7A97: d <= 8'h41;
                15'h7A98: d <= 8'h49; 15'h7A99: d <= 8'h4D; 15'h7A9A: d <= 8'h42; 15'h7A9B: d <= 8'h46;
                15'h7A9C: d <= 8'h4E; 15'h7A9D: d <= 8'h43; 15'h7A9E: d <= 8'h47; 15'h7A9F: d <= 8'h4B;
                15'h7AA0: d <= 8'h50; 15'h7AA1: d <= 8'h55; 15'h7AA2: d <= 8'h5A; 15'h7AA3: d <= 8'h5F;
                15'h7AA4: d <= 8'h60; 15'h7AA5: d <= 8'h65; 15'h7AA6: d <= 8'h6A; 15'h7AA7: d <= 8'h6F;
                15'h7AA8: d <= 8'h74; 15'h7AA9: d <= 8'h78; 15'h7AAA: d <= 8'h7C; 15'h7AAB: d <= 8'h71;
                15'h7AAC: d <= 8'h79; 15'h7AAD: d <= 8'h7D; 15'h7AAE: d <= 8'h72; 15'h7AAF: d <= 8'h76;
                15'h7AB0: d <= 8'h7E; 15'h7AB1: d <= 8'h73; 15'h7AB2: d <= 8'h77; 15'h7AB3: d <= 8'h7B;
                15'h7AB4: d <= 8'h84; 15'h7AB5: d <= 8'h88; 15'h7AB6: d <= 8'h8C; 15'h7AB7: d <= 8'h81;
                15'h7AB8: d <= 8'h89; 15'h7AB9: d <= 8'h8D; 15'h7ABA: d <= 8'h82; 15'h7ABB: d <= 8'h86;
                15'h7ABC: d <= 8'h8E; 15'h7ABD: d <= 8'h83; 15'h7ABE: d <= 8'h87; 15'h7ABF: d <= 8'h8B;
                15'h7AC0: d <= 8'h90; 15'h7AC1: d <= 8'h95; 15'h7AC2: d <= 8'h9A; 15'h7AC3: d <= 8'h9F;
                15'h7AC4: d <= 8'hA4; 15'h7AC5: d <= 8'hA8; 15'h7AC6: d <= 8'hAC; 15'h7AC7: d <= 8'hA1;
                15'h7AC8: d <= 8'hA9; 15'h7AC9: d <= 8'hAD; 15'h7ACA: d <= 8'hA2; 15'h7ACB: d <= 8'hA6;
                15'h7ACC: d <= 8'hAE; 15'h7ACD: d <= 8'hA3; 15'h7ACE: d <= 8'hA7; 15'h7ACF: d <= 8'hAB;
                15'h7AD0: d <= 8'hB4; 15'h7AD1: d <= 8'hB8; 15'h7AD2: d <= 8'hBC; 15'h7AD3: d <= 8'hB1;
                15'h7AD4: d <= 8'hB9; 15'h7AD5: d <= 8'hBD; 15'h7AD6: d <= 8'hB2; 15'h7AD7: d <= 8'hB6;
                15'h7AD8: d <= 8'hBE; 15'h7AD9: d <= 8'hB3; 15'h7ADA: d <= 8'hB7; 15'h7ADB: d <= 8'hBB;
                15'h7ADC: d <= 8'hC4; 15'h7ADD: d <= 8'hC8; 15'h7ADE: d <= 8'hCC; 15'h7ADF: d <= 8'hC1;
                15'h7AE0: d <= 8'hC9; 15'h7AE1: d <= 8'hCD; 15'h7AE2: d <= 8'hC2; 15'h7AE3: d <= 8'hC6;
                15'h7AE4: d <= 8'hCE; 15'h7AE5: d <= 8'hC3; 15'h7AE6: d <= 8'hC7; 15'h7AE7: d <= 8'hCB;
                15'h7AE8: d <= 8'hC0; 15'h7AE9: d <= 8'hC5; 15'h7AEA: d <= 8'hCA; 15'h7AEB: d <= 8'hCF;
                15'h7AEC: d <= 8'hD0; 15'h7AED: d <= 8'hD5; 15'h7AEE: d <= 8'hDA; 15'h7AEF: d <= 8'hDF;
                15'h7AF0: d <= 8'h74; 15'h7AF1: d <= 8'h78; 15'h7AF2: d <= 8'h7C; 15'h7AF3: d <= 8'h71;
                15'h7AF4: d <= 8'h79; 15'h7AF5: d <= 8'h7D; 15'h7AF6: d <= 8'h72; 15'h7AF7: d <= 8'h76;
                15'h7AF8: d <= 8'h7E; 15'h7AF9: d <= 8'h73; 15'h7AFA: d <= 8'h77; 15'h7AFB: d <= 8'h7B;
                15'h7AFC: d <= 8'hA0; 15'h7AFD: d <= 8'hA5; 15'h7AFE: d <= 8'hAA; 15'h7AFF: d <= 8'hAF;
                15'h7B00: d <= 8'h00; 15'h7B01: d <= 8'h00; 15'h7B02: d <= 8'h00; 15'h7B03: d <= 8'h00;
                15'h7B04: d <= 8'h00; 15'h7B05: d <= 8'h00; 15'h7B06: d <= 8'h00; 15'h7B07: d <= 8'h00;
                15'h7B08: d <= 8'h00; 15'h7B09: d <= 8'h00; 15'h7B0A: d <= 8'h00; 15'h7B0B: d <= 8'h00;
                15'h7B0C: d <= 8'h00; 15'h7B0D: d <= 8'h00; 15'h7B0E: d <= 8'h00; 15'h7B0F: d <= 8'h00;
                15'h7B10: d <= 8'h00; 15'h7B11: d <= 8'h00; 15'h7B12: d <= 8'h00; 15'h7B13: d <= 8'h00;
                15'h7B14: d <= 8'h00; 15'h7B15: d <= 8'h00; 15'h7B16: d <= 8'h00; 15'h7B17: d <= 8'h00;
                15'h7B18: d <= 8'h00; 15'h7B19: d <= 8'h00; 15'h7B1A: d <= 8'h00; 15'h7B1B: d <= 8'h00;
                15'h7B1C: d <= 8'h00; 15'h7B1D: d <= 8'h00; 15'h7B1E: d <= 8'h00; 15'h7B1F: d <= 8'h00;
                15'h7B20: d <= 8'h00; 15'h7B21: d <= 8'h00; 15'h7B22: d <= 8'h00; 15'h7B23: d <= 8'h00;
                15'h7B24: d <= 8'h00; 15'h7B25: d <= 8'h00; 15'h7B26: d <= 8'h00; 15'h7B27: d <= 8'h00;
                15'h7B28: d <= 8'h00; 15'h7B29: d <= 8'h00; 15'h7B2A: d <= 8'h00; 15'h7B2B: d <= 8'h00;
                15'h7B2C: d <= 8'h00; 15'h7B2D: d <= 8'h00; 15'h7B2E: d <= 8'h00; 15'h7B2F: d <= 8'h7B;
                15'h7B30: d <= 8'h00; 15'h7B31: d <= 8'h00; 15'h7B32: d <= 8'h00; 15'h7B33: d <= 8'h00;
                15'h7B34: d <= 8'h00; 15'h7B35: d <= 8'h00; 15'h7B36: d <= 8'h00; 15'h7B37: d <= 8'h00;
                15'h7B38: d <= 8'h00; 15'h7B39: d <= 8'h00; 15'h7B3A: d <= 8'h00; 15'h7B3B: d <= 8'h00;
                15'h7B3C: d <= 8'h00; 15'h7B3D: d <= 8'h00; 15'h7B3E: d <= 8'h00; 15'h7B3F: d <= 8'h00;
                15'h7B40: d <= 8'h00; 15'h7B41: d <= 8'h00; 15'h7B42: d <= 8'h00; 15'h7B43: d <= 8'h00;
                15'h7B44: d <= 8'h00; 15'h7B45: d <= 8'h00; 15'h7B46: d <= 8'h00; 15'h7B47: d <= 8'h00;
                15'h7B48: d <= 8'h00; 15'h7B49: d <= 8'h00; 15'h7B4A: d <= 8'h00; 15'h7B4B: d <= 8'h00;
                15'h7B4C: d <= 8'h00; 15'h7B4D: d <= 8'h00; 15'h7B4E: d <= 8'h00; 15'h7B4F: d <= 8'h00;
                15'h7B50: d <= 8'h00; 15'h7B51: d <= 8'h00; 15'h7B52: d <= 8'h00; 15'h7B53: d <= 8'h00;
                15'h7B54: d <= 8'h00; 15'h7B55: d <= 8'h00; 15'h7B56: d <= 8'h00; 15'h7B57: d <= 8'h00;
                15'h7B58: d <= 8'h45; 15'h7B59: d <= 8'h35; 15'h7B5A: d <= 8'h32; 15'h7B5B: d <= 8'h00;
                15'h7B5C: d <= 8'h00; 15'h7B5D: d <= 8'h00; 15'h7B5E: d <= 8'h00; 15'h7B5F: d <= 8'h00;
                15'h7B60: d <= 8'h00; 15'h7B61: d <= 8'h00; 15'h7B62: d <= 8'h00; 15'h7B63: d <= 8'h00;
                15'h7B64: d <= 8'h00; 15'h7B65: d <= 8'h00; 15'h7B66: d <= 8'h00; 15'h7B67: d <= 8'h00;
                15'h7B68: d <= 8'h00; 15'h7B69: d <= 8'h00; 15'h7B6A: d <= 8'h00; 15'h7B6B: d <= 8'h00;
                15'h7B6C: d <= 8'h00; 15'h7B6D: d <= 8'h00; 15'h7B6E: d <= 8'h00; 15'h7B6F: d <= 8'h00;
                15'h7B70: d <= 8'h00; 15'h7B71: d <= 8'h00; 15'h7B72: d <= 8'h00; 15'h7B73: d <= 8'h00;
                15'h7B74: d <= 8'h00; 15'h7B75: d <= 8'h00; 15'h7B76: d <= 8'h00; 15'h7B77: d <= 8'h00;
                15'h7B78: d <= 8'h00; 15'h7B79: d <= 8'h00; 15'h7B7A: d <= 8'h00; 15'h7B7B: d <= 8'h00;
                15'h7B7C: d <= 8'h00; 15'h7B7D: d <= 8'h00; 15'h7B7E: d <= 8'h00; 15'h7B7F: d <= 8'hE0;
                15'h7B80: d <= 8'h10; 15'h7B81: d <= 8'h15; 15'h7B82: d <= 8'h1A; 15'h7B83: d <= 8'h1F;
                15'h7B84: d <= 8'h20; 15'h7B85: d <= 8'h25; 15'h7B86: d <= 8'h2A; 15'h7B87: d <= 8'h2F;
                15'h7B88: d <= 8'h34; 15'h7B89: d <= 8'h38; 15'h7B8A: d <= 8'h3C; 15'h7B8B: d <= 8'h31;
                15'h7B8C: d <= 8'h39; 15'h7B8D: d <= 8'h3D; 15'h7B8E: d <= 8'h32; 15'h7B8F: d <= 8'h36;
                15'h7B90: d <= 8'h3E; 15'h7B91: d <= 8'h33; 15'h7B92: d <= 8'h37; 15'h7B93: d <= 8'h3B;
                15'h7B94: d <= 8'h44; 15'h7B95: d <= 8'h48; 15'h7B96: d <= 8'h4C; 15'h7B97: d <= 8'h41;
                15'h7B98: d <= 8'h49; 15'h7B99: d <= 8'h4D; 15'h7B9A: d <= 8'h42; 15'h7B9B: d <= 8'h46;
                15'h7B9C: d <= 8'h4E; 15'h7B9D: d <= 8'h43; 15'h7B9E: d <= 8'h47; 15'h7B9F: d <= 8'h4B;
                15'h7BA0: d <= 8'h50; 15'h7BA1: d <= 8'h55; 15'h7BA2: d <= 8'h5A; 15'h7BA3: d <= 8'h5F;
                15'h7BA4: d <= 8'h60; 15'h7BA5: d <= 8'h65; 15'h7BA6: d <= 8'h6A; 15'h7BA7: d <= 8'h6F;
                15'h7BA8: d <= 8'h74; 15'h7BA9: d <= 8'h78; 15'h7BAA: d <= 8'h7C; 15'h7BAB: d <= 8'h71;
                15'h7BAC: d <= 8'h79; 15'h7BAD: d <= 8'h7D; 15'h7BAE: d <= 8'h72; 15'h7BAF: d <= 8'h76;
                15'h7BB0: d <= 8'h7E; 15'h7BB1: d <= 8'h73; 15'h7BB2: d <= 8'h77; 15'h7BB3: d <= 8'h7B;
                15'h7BB4: d <= 8'h84; 15'h7BB5: d <= 8'h88; 15'h7BB6: d <= 8'h8C; 15'h7BB7: d <= 8'h81;
                15'h7BB8: d <= 8'h89; 15'h7BB9: d <= 8'h8D; 15'h7BBA: d <= 8'h82; 15'h7BBB: d <= 8'h86;
                15'h7BBC: d <= 8'h8E; 15'h7BBD: d <= 8'h83; 15'h7BBE: d <= 8'h87; 15'h7BBF: d <= 8'h8B;
                15'h7BC0: d <= 8'h90; 15'h7BC1: d <= 8'h95; 15'h7BC2: d <= 8'h9A; 15'h7BC3: d <= 8'h9F;
                15'h7BC4: d <= 8'hA4; 15'h7BC5: d <= 8'hA8; 15'h7BC6: d <= 8'hAC; 15'h7BC7: d <= 8'hA1;
                15'h7BC8: d <= 8'hA9; 15'h7BC9: d <= 8'hAD; 15'h7BCA: d <= 8'hA2; 15'h7BCB: d <= 8'hA6;
                15'h7BCC: d <= 8'hAE; 15'h7BCD: d <= 8'hA3; 15'h7BCE: d <= 8'hA7; 15'h7BCF: d <= 8'hAB;
                15'h7BD0: d <= 8'hB4; 15'h7BD1: d <= 8'hB8; 15'h7BD2: d <= 8'hBC; 15'h7BD3: d <= 8'hB1;
                15'h7BD4: d <= 8'hB9; 15'h7BD5: d <= 8'hBD; 15'h7BD6: d <= 8'hB2; 15'h7BD7: d <= 8'hB6;
                15'h7BD8: d <= 8'hBE; 15'h7BD9: d <= 8'hB3; 15'h7BDA: d <= 8'hB7; 15'h7BDB: d <= 8'hBB;
                15'h7BDC: d <= 8'hC4; 15'h7BDD: d <= 8'hC8; 15'h7BDE: d <= 8'hCC; 15'h7BDF: d <= 8'hC1;
                15'h7BE0: d <= 8'hC9; 15'h7BE1: d <= 8'hCD; 15'h7BE2: d <= 8'hC2; 15'h7BE3: d <= 8'hC6;
                15'h7BE4: d <= 8'hCE; 15'h7BE5: d <= 8'hC3; 15'h7BE6: d <= 8'hC7; 15'h7BE7: d <= 8'hCB;
                15'h7BE8: d <= 8'hC0; 15'h7BE9: d <= 8'hC5; 15'h7BEA: d <= 8'hCA; 15'h7BEB: d <= 8'hCF;
                15'h7BEC: d <= 8'hD0; 15'h7BED: d <= 8'hD5; 15'h7BEE: d <= 8'hDA; 15'h7BEF: d <= 8'hDF;
                15'h7BF0: d <= 8'h74; 15'h7BF1: d <= 8'h78; 15'h7BF2: d <= 8'h7C; 15'h7BF3: d <= 8'h71;
                15'h7BF4: d <= 8'h79; 15'h7BF5: d <= 8'h7D; 15'h7BF6: d <= 8'h72; 15'h7BF7: d <= 8'h76;
                15'h7BF8: d <= 8'h7E; 15'h7BF9: d <= 8'h73; 15'h7BFA: d <= 8'h77; 15'h7BFB: d <= 8'h7B;
                15'h7BFC: d <= 8'hA0; 15'h7BFD: d <= 8'hA5; 15'h7BFE: d <= 8'hAA; 15'h7BFF: d <= 8'hAF;
                15'h7C00: d <= 8'h00; 15'h7C01: d <= 8'h00; 15'h7C02: d <= 8'h00; 15'h7C03: d <= 8'h00;
                15'h7C04: d <= 8'h00; 15'h7C05: d <= 8'h00; 15'h7C06: d <= 8'h00; 15'h7C07: d <= 8'h00;
                15'h7C08: d <= 8'h00; 15'h7C09: d <= 8'h00; 15'h7C0A: d <= 8'h00; 15'h7C0B: d <= 8'h00;
                15'h7C0C: d <= 8'h00; 15'h7C0D: d <= 8'h00; 15'h7C0E: d <= 8'h00; 15'h7C0F: d <= 8'h00;
                15'h7C10: d <= 8'h00; 15'h7C11: d <= 8'h00; 15'h7C12: d <= 8'h00; 15'h7C13: d <= 8'h00;
                15'h7C14: d <= 8'h00; 15'h7C15: d <= 8'h00; 15'h7C16: d <= 8'h00; 15'h7C17: d <= 8'h00;
                15'h7C18: d <= 8'h00; 15'h7C19: d <= 8'h00; 15'h7C1A: d <= 8'h00; 15'h7C1B: d <= 8'h00;
                15'h7C1C: d <= 8'h00; 15'h7C1D: d <= 8'h00; 15'h7C1E: d <= 8'h00; 15'h7C1F: d <= 8'h00;
                15'h7C20: d <= 8'h00; 15'h7C21: d <= 8'h00; 15'h7C22: d <= 8'h00; 15'h7C23: d <= 8'h00;
                15'h7C24: d <= 8'h00; 15'h7C25: d <= 8'h00; 15'h7C26: d <= 8'h00; 15'h7C27: d <= 8'h00;
                15'h7C28: d <= 8'h00; 15'h7C29: d <= 8'h00; 15'h7C2A: d <= 8'h00; 15'h7C2B: d <= 8'h00;
                15'h7C2C: d <= 8'h00; 15'h7C2D: d <= 8'h00; 15'h7C2E: d <= 8'h00; 15'h7C2F: d <= 8'h7B;
                15'h7C30: d <= 8'h00; 15'h7C31: d <= 8'h00; 15'h7C32: d <= 8'h00; 15'h7C33: d <= 8'h00;
                15'h7C34: d <= 8'h00; 15'h7C35: d <= 8'h00; 15'h7C36: d <= 8'h00; 15'h7C37: d <= 8'h00;
                15'h7C38: d <= 8'h00; 15'h7C39: d <= 8'h00; 15'h7C3A: d <= 8'h00; 15'h7C3B: d <= 8'h00;
                15'h7C3C: d <= 8'h00; 15'h7C3D: d <= 8'h00; 15'h7C3E: d <= 8'h00; 15'h7C3F: d <= 8'h00;
                15'h7C40: d <= 8'h00; 15'h7C41: d <= 8'h00; 15'h7C42: d <= 8'h00; 15'h7C43: d <= 8'h00;
                15'h7C44: d <= 8'h00; 15'h7C45: d <= 8'h00; 15'h7C46: d <= 8'h00; 15'h7C47: d <= 8'h00;
                15'h7C48: d <= 8'h00; 15'h7C49: d <= 8'h00; 15'h7C4A: d <= 8'h00; 15'h7C4B: d <= 8'h00;
                15'h7C4C: d <= 8'h00; 15'h7C4D: d <= 8'h00; 15'h7C4E: d <= 8'h00; 15'h7C4F: d <= 8'h00;
                15'h7C50: d <= 8'h00; 15'h7C51: d <= 8'h00; 15'h7C52: d <= 8'h00; 15'h7C53: d <= 8'h00;
                15'h7C54: d <= 8'h00; 15'h7C55: d <= 8'h00; 15'h7C56: d <= 8'h00; 15'h7C57: d <= 8'h00;
                15'h7C58: d <= 8'h45; 15'h7C59: d <= 8'h35; 15'h7C5A: d <= 8'h32; 15'h7C5B: d <= 8'h00;
                15'h7C5C: d <= 8'h00; 15'h7C5D: d <= 8'h00; 15'h7C5E: d <= 8'h00; 15'h7C5F: d <= 8'h00;
                15'h7C60: d <= 8'h00; 15'h7C61: d <= 8'h00; 15'h7C62: d <= 8'h00; 15'h7C63: d <= 8'h00;
                15'h7C64: d <= 8'h00; 15'h7C65: d <= 8'h00; 15'h7C66: d <= 8'h00; 15'h7C67: d <= 8'h00;
                15'h7C68: d <= 8'h00; 15'h7C69: d <= 8'h00; 15'h7C6A: d <= 8'h00; 15'h7C6B: d <= 8'h00;
                15'h7C6C: d <= 8'h00; 15'h7C6D: d <= 8'h00; 15'h7C6E: d <= 8'h00; 15'h7C6F: d <= 8'h00;
                15'h7C70: d <= 8'h00; 15'h7C71: d <= 8'h00; 15'h7C72: d <= 8'h00; 15'h7C73: d <= 8'h00;
                15'h7C74: d <= 8'h00; 15'h7C75: d <= 8'h00; 15'h7C76: d <= 8'h00; 15'h7C77: d <= 8'h00;
                15'h7C78: d <= 8'h00; 15'h7C79: d <= 8'h00; 15'h7C7A: d <= 8'h00; 15'h7C7B: d <= 8'h00;
                15'h7C7C: d <= 8'h00; 15'h7C7D: d <= 8'h00; 15'h7C7E: d <= 8'h00; 15'h7C7F: d <= 8'hE0;
                15'h7C80: d <= 8'h10; 15'h7C81: d <= 8'h15; 15'h7C82: d <= 8'h1A; 15'h7C83: d <= 8'h1F;
                15'h7C84: d <= 8'h20; 15'h7C85: d <= 8'h25; 15'h7C86: d <= 8'h2A; 15'h7C87: d <= 8'h2F;
                15'h7C88: d <= 8'h34; 15'h7C89: d <= 8'h38; 15'h7C8A: d <= 8'h3C; 15'h7C8B: d <= 8'h31;
                15'h7C8C: d <= 8'h39; 15'h7C8D: d <= 8'h3D; 15'h7C8E: d <= 8'h32; 15'h7C8F: d <= 8'h36;
                15'h7C90: d <= 8'h3E; 15'h7C91: d <= 8'h33; 15'h7C92: d <= 8'h37; 15'h7C93: d <= 8'h3B;
                15'h7C94: d <= 8'h44; 15'h7C95: d <= 8'h48; 15'h7C96: d <= 8'h4C; 15'h7C97: d <= 8'h41;
                15'h7C98: d <= 8'h49; 15'h7C99: d <= 8'h4D; 15'h7C9A: d <= 8'h42; 15'h7C9B: d <= 8'h46;
                15'h7C9C: d <= 8'h4E; 15'h7C9D: d <= 8'h43; 15'h7C9E: d <= 8'h47; 15'h7C9F: d <= 8'h4B;
                15'h7CA0: d <= 8'h50; 15'h7CA1: d <= 8'h55; 15'h7CA2: d <= 8'h5A; 15'h7CA3: d <= 8'h5F;
                15'h7CA4: d <= 8'h60; 15'h7CA5: d <= 8'h65; 15'h7CA6: d <= 8'h6A; 15'h7CA7: d <= 8'h6F;
                15'h7CA8: d <= 8'h74; 15'h7CA9: d <= 8'h78; 15'h7CAA: d <= 8'h7C; 15'h7CAB: d <= 8'h71;
                15'h7CAC: d <= 8'h79; 15'h7CAD: d <= 8'h7D; 15'h7CAE: d <= 8'h72; 15'h7CAF: d <= 8'h76;
                15'h7CB0: d <= 8'h7E; 15'h7CB1: d <= 8'h73; 15'h7CB2: d <= 8'h77; 15'h7CB3: d <= 8'h7B;
                15'h7CB4: d <= 8'h84; 15'h7CB5: d <= 8'h88; 15'h7CB6: d <= 8'h8C; 15'h7CB7: d <= 8'h81;
                15'h7CB8: d <= 8'h89; 15'h7CB9: d <= 8'h8D; 15'h7CBA: d <= 8'h82; 15'h7CBB: d <= 8'h86;
                15'h7CBC: d <= 8'h8E; 15'h7CBD: d <= 8'h83; 15'h7CBE: d <= 8'h87; 15'h7CBF: d <= 8'h8B;
                15'h7CC0: d <= 8'h90; 15'h7CC1: d <= 8'h95; 15'h7CC2: d <= 8'h9A; 15'h7CC3: d <= 8'h9F;
                15'h7CC4: d <= 8'hA4; 15'h7CC5: d <= 8'hA8; 15'h7CC6: d <= 8'hAC; 15'h7CC7: d <= 8'hA1;
                15'h7CC8: d <= 8'hA9; 15'h7CC9: d <= 8'hAD; 15'h7CCA: d <= 8'hA2; 15'h7CCB: d <= 8'hA6;
                15'h7CCC: d <= 8'hAE; 15'h7CCD: d <= 8'hA3; 15'h7CCE: d <= 8'hA7; 15'h7CCF: d <= 8'hAB;
                15'h7CD0: d <= 8'hB4; 15'h7CD1: d <= 8'hB8; 15'h7CD2: d <= 8'hBC; 15'h7CD3: d <= 8'hB1;
                15'h7CD4: d <= 8'hB9; 15'h7CD5: d <= 8'hBD; 15'h7CD6: d <= 8'hB2; 15'h7CD7: d <= 8'hB6;
                15'h7CD8: d <= 8'hBE; 15'h7CD9: d <= 8'hB3; 15'h7CDA: d <= 8'hB7; 15'h7CDB: d <= 8'hBB;
                15'h7CDC: d <= 8'hC4; 15'h7CDD: d <= 8'hC8; 15'h7CDE: d <= 8'hCC; 15'h7CDF: d <= 8'hC1;
                15'h7CE0: d <= 8'hC9; 15'h7CE1: d <= 8'hCD; 15'h7CE2: d <= 8'hC2; 15'h7CE3: d <= 8'hC6;
                15'h7CE4: d <= 8'hCE; 15'h7CE5: d <= 8'hC3; 15'h7CE6: d <= 8'hC7; 15'h7CE7: d <= 8'hCB;
                15'h7CE8: d <= 8'hC0; 15'h7CE9: d <= 8'hC5; 15'h7CEA: d <= 8'hCA; 15'h7CEB: d <= 8'hCF;
                15'h7CEC: d <= 8'hD0; 15'h7CED: d <= 8'hD5; 15'h7CEE: d <= 8'hDA; 15'h7CEF: d <= 8'hDF;
                15'h7CF0: d <= 8'h74; 15'h7CF1: d <= 8'h78; 15'h7CF2: d <= 8'h7C; 15'h7CF3: d <= 8'h71;
                15'h7CF4: d <= 8'h79; 15'h7CF5: d <= 8'h7D; 15'h7CF6: d <= 8'h72; 15'h7CF7: d <= 8'h76;
                15'h7CF8: d <= 8'h7E; 15'h7CF9: d <= 8'h73; 15'h7CFA: d <= 8'h77; 15'h7CFB: d <= 8'h7B;
                15'h7CFC: d <= 8'hA0; 15'h7CFD: d <= 8'hA5; 15'h7CFE: d <= 8'hAA; 15'h7CFF: d <= 8'hAF;
                15'h7D00: d <= 8'h00; 15'h7D01: d <= 8'h00; 15'h7D02: d <= 8'h00; 15'h7D03: d <= 8'h00;
                15'h7D04: d <= 8'h00; 15'h7D05: d <= 8'h00; 15'h7D06: d <= 8'h00; 15'h7D07: d <= 8'h00;
                15'h7D08: d <= 8'h00; 15'h7D09: d <= 8'h00; 15'h7D0A: d <= 8'h00; 15'h7D0B: d <= 8'h00;
                15'h7D0C: d <= 8'h00; 15'h7D0D: d <= 8'h00; 15'h7D0E: d <= 8'h00; 15'h7D0F: d <= 8'h00;
                15'h7D10: d <= 8'h00; 15'h7D11: d <= 8'h00; 15'h7D12: d <= 8'h00; 15'h7D13: d <= 8'h00;
                15'h7D14: d <= 8'h00; 15'h7D15: d <= 8'h00; 15'h7D16: d <= 8'h00; 15'h7D17: d <= 8'h00;
                15'h7D18: d <= 8'h00; 15'h7D19: d <= 8'h00; 15'h7D1A: d <= 8'h00; 15'h7D1B: d <= 8'h00;
                15'h7D1C: d <= 8'h00; 15'h7D1D: d <= 8'h00; 15'h7D1E: d <= 8'h00; 15'h7D1F: d <= 8'h00;
                15'h7D20: d <= 8'h00; 15'h7D21: d <= 8'h00; 15'h7D22: d <= 8'h00; 15'h7D23: d <= 8'h00;
                15'h7D24: d <= 8'h00; 15'h7D25: d <= 8'h00; 15'h7D26: d <= 8'h00; 15'h7D27: d <= 8'h00;
                15'h7D28: d <= 8'h00; 15'h7D29: d <= 8'h00; 15'h7D2A: d <= 8'h00; 15'h7D2B: d <= 8'h00;
                15'h7D2C: d <= 8'h00; 15'h7D2D: d <= 8'h00; 15'h7D2E: d <= 8'h00; 15'h7D2F: d <= 8'h7B;
                15'h7D30: d <= 8'h00; 15'h7D31: d <= 8'h00; 15'h7D32: d <= 8'h00; 15'h7D33: d <= 8'h00;
                15'h7D34: d <= 8'h00; 15'h7D35: d <= 8'h00; 15'h7D36: d <= 8'h00; 15'h7D37: d <= 8'h00;
                15'h7D38: d <= 8'h00; 15'h7D39: d <= 8'h00; 15'h7D3A: d <= 8'h00; 15'h7D3B: d <= 8'h00;
                15'h7D3C: d <= 8'h00; 15'h7D3D: d <= 8'h00; 15'h7D3E: d <= 8'h00; 15'h7D3F: d <= 8'h00;
                15'h7D40: d <= 8'h00; 15'h7D41: d <= 8'h00; 15'h7D42: d <= 8'h00; 15'h7D43: d <= 8'h00;
                15'h7D44: d <= 8'h00; 15'h7D45: d <= 8'h00; 15'h7D46: d <= 8'h00; 15'h7D47: d <= 8'h00;
                15'h7D48: d <= 8'h00; 15'h7D49: d <= 8'h00; 15'h7D4A: d <= 8'h00; 15'h7D4B: d <= 8'h00;
                15'h7D4C: d <= 8'h00; 15'h7D4D: d <= 8'h00; 15'h7D4E: d <= 8'h00; 15'h7D4F: d <= 8'h00;
                15'h7D50: d <= 8'h00; 15'h7D51: d <= 8'h00; 15'h7D52: d <= 8'h00; 15'h7D53: d <= 8'h00;
                15'h7D54: d <= 8'h00; 15'h7D55: d <= 8'h00; 15'h7D56: d <= 8'h00; 15'h7D57: d <= 8'h00;
                15'h7D58: d <= 8'h45; 15'h7D59: d <= 8'h35; 15'h7D5A: d <= 8'h32; 15'h7D5B: d <= 8'h00;
                15'h7D5C: d <= 8'h00; 15'h7D5D: d <= 8'h00; 15'h7D5E: d <= 8'h00; 15'h7D5F: d <= 8'h00;
                15'h7D60: d <= 8'h00; 15'h7D61: d <= 8'h00; 15'h7D62: d <= 8'h00; 15'h7D63: d <= 8'h00;
                15'h7D64: d <= 8'h00; 15'h7D65: d <= 8'h00; 15'h7D66: d <= 8'h00; 15'h7D67: d <= 8'h00;
                15'h7D68: d <= 8'h00; 15'h7D69: d <= 8'h00; 15'h7D6A: d <= 8'h00; 15'h7D6B: d <= 8'h00;
                15'h7D6C: d <= 8'h00; 15'h7D6D: d <= 8'h00; 15'h7D6E: d <= 8'h00; 15'h7D6F: d <= 8'h00;
                15'h7D70: d <= 8'h00; 15'h7D71: d <= 8'h00; 15'h7D72: d <= 8'h00; 15'h7D73: d <= 8'h00;
                15'h7D74: d <= 8'h00; 15'h7D75: d <= 8'h00; 15'h7D76: d <= 8'h00; 15'h7D77: d <= 8'h00;
                15'h7D78: d <= 8'h00; 15'h7D79: d <= 8'h00; 15'h7D7A: d <= 8'h00; 15'h7D7B: d <= 8'h00;
                15'h7D7C: d <= 8'h00; 15'h7D7D: d <= 8'h00; 15'h7D7E: d <= 8'h00; 15'h7D7F: d <= 8'hE0;
                15'h7D80: d <= 8'h10; 15'h7D81: d <= 8'h15; 15'h7D82: d <= 8'h1A; 15'h7D83: d <= 8'h1F;
                15'h7D84: d <= 8'h20; 15'h7D85: d <= 8'h25; 15'h7D86: d <= 8'h2A; 15'h7D87: d <= 8'h2F;
                15'h7D88: d <= 8'h34; 15'h7D89: d <= 8'h38; 15'h7D8A: d <= 8'h3C; 15'h7D8B: d <= 8'h31;
                15'h7D8C: d <= 8'h39; 15'h7D8D: d <= 8'h3D; 15'h7D8E: d <= 8'h32; 15'h7D8F: d <= 8'h36;
                15'h7D90: d <= 8'h3E; 15'h7D91: d <= 8'h33; 15'h7D92: d <= 8'h37; 15'h7D93: d <= 8'h3B;
                15'h7D94: d <= 8'h44; 15'h7D95: d <= 8'h48; 15'h7D96: d <= 8'h4C; 15'h7D97: d <= 8'h41;
                15'h7D98: d <= 8'h49; 15'h7D99: d <= 8'h4D; 15'h7D9A: d <= 8'h42; 15'h7D9B: d <= 8'h46;
                15'h7D9C: d <= 8'h4E; 15'h7D9D: d <= 8'h43; 15'h7D9E: d <= 8'h47; 15'h7D9F: d <= 8'h4B;
                15'h7DA0: d <= 8'h50; 15'h7DA1: d <= 8'h55; 15'h7DA2: d <= 8'h5A; 15'h7DA3: d <= 8'h5F;
                15'h7DA4: d <= 8'h60; 15'h7DA5: d <= 8'h65; 15'h7DA6: d <= 8'h6A; 15'h7DA7: d <= 8'h6F;
                15'h7DA8: d <= 8'h74; 15'h7DA9: d <= 8'h78; 15'h7DAA: d <= 8'h7C; 15'h7DAB: d <= 8'h71;
                15'h7DAC: d <= 8'h79; 15'h7DAD: d <= 8'h7D; 15'h7DAE: d <= 8'h72; 15'h7DAF: d <= 8'h76;
                15'h7DB0: d <= 8'h7E; 15'h7DB1: d <= 8'h73; 15'h7DB2: d <= 8'h77; 15'h7DB3: d <= 8'h7B;
                15'h7DB4: d <= 8'h84; 15'h7DB5: d <= 8'h88; 15'h7DB6: d <= 8'h8C; 15'h7DB7: d <= 8'h81;
                15'h7DB8: d <= 8'h89; 15'h7DB9: d <= 8'h8D; 15'h7DBA: d <= 8'h82; 15'h7DBB: d <= 8'h86;
                15'h7DBC: d <= 8'h8E; 15'h7DBD: d <= 8'h83; 15'h7DBE: d <= 8'h87; 15'h7DBF: d <= 8'h8B;
                15'h7DC0: d <= 8'h90; 15'h7DC1: d <= 8'h95; 15'h7DC2: d <= 8'h9A; 15'h7DC3: d <= 8'h9F;
                15'h7DC4: d <= 8'hA4; 15'h7DC5: d <= 8'hA8; 15'h7DC6: d <= 8'hAC; 15'h7DC7: d <= 8'hA1;
                15'h7DC8: d <= 8'hA9; 15'h7DC9: d <= 8'hAD; 15'h7DCA: d <= 8'hA2; 15'h7DCB: d <= 8'hA6;
                15'h7DCC: d <= 8'hAE; 15'h7DCD: d <= 8'hA3; 15'h7DCE: d <= 8'hA7; 15'h7DCF: d <= 8'hAB;
                15'h7DD0: d <= 8'hB4; 15'h7DD1: d <= 8'hB8; 15'h7DD2: d <= 8'hBC; 15'h7DD3: d <= 8'hB1;
                15'h7DD4: d <= 8'hB9; 15'h7DD5: d <= 8'hBD; 15'h7DD6: d <= 8'hB2; 15'h7DD7: d <= 8'hB6;
                15'h7DD8: d <= 8'hBE; 15'h7DD9: d <= 8'hB3; 15'h7DDA: d <= 8'hB7; 15'h7DDB: d <= 8'hBB;
                15'h7DDC: d <= 8'hC4; 15'h7DDD: d <= 8'hC8; 15'h7DDE: d <= 8'hCC; 15'h7DDF: d <= 8'hC1;
                15'h7DE0: d <= 8'hC9; 15'h7DE1: d <= 8'hCD; 15'h7DE2: d <= 8'hC2; 15'h7DE3: d <= 8'hC6;
                15'h7DE4: d <= 8'hCE; 15'h7DE5: d <= 8'hC3; 15'h7DE6: d <= 8'hC7; 15'h7DE7: d <= 8'hCB;
                15'h7DE8: d <= 8'hC0; 15'h7DE9: d <= 8'hC5; 15'h7DEA: d <= 8'hCA; 15'h7DEB: d <= 8'hCF;
                15'h7DEC: d <= 8'hD0; 15'h7DED: d <= 8'hD5; 15'h7DEE: d <= 8'hDA; 15'h7DEF: d <= 8'hDF;
                15'h7DF0: d <= 8'h74; 15'h7DF1: d <= 8'h78; 15'h7DF2: d <= 8'h7C; 15'h7DF3: d <= 8'h71;
                15'h7DF4: d <= 8'h79; 15'h7DF5: d <= 8'h7D; 15'h7DF6: d <= 8'h72; 15'h7DF7: d <= 8'h76;
                15'h7DF8: d <= 8'h7E; 15'h7DF9: d <= 8'h73; 15'h7DFA: d <= 8'h77; 15'h7DFB: d <= 8'h7B;
                15'h7DFC: d <= 8'hA0; 15'h7DFD: d <= 8'hA5; 15'h7DFE: d <= 8'hAA; 15'h7DFF: d <= 8'hAF;
                15'h7E00: d <= 8'h00; 15'h7E01: d <= 8'h00; 15'h7E02: d <= 8'h00; 15'h7E03: d <= 8'h00;
                15'h7E04: d <= 8'h00; 15'h7E05: d <= 8'h00; 15'h7E06: d <= 8'h00; 15'h7E07: d <= 8'h00;
                15'h7E08: d <= 8'h00; 15'h7E09: d <= 8'h00; 15'h7E0A: d <= 8'h00; 15'h7E0B: d <= 8'h00;
                15'h7E0C: d <= 8'h00; 15'h7E0D: d <= 8'h00; 15'h7E0E: d <= 8'h00; 15'h7E0F: d <= 8'h00;
                15'h7E10: d <= 8'h00; 15'h7E11: d <= 8'h00; 15'h7E12: d <= 8'h00; 15'h7E13: d <= 8'h00;
                15'h7E14: d <= 8'h00; 15'h7E15: d <= 8'h00; 15'h7E16: d <= 8'h00; 15'h7E17: d <= 8'h00;
                15'h7E18: d <= 8'h00; 15'h7E19: d <= 8'h00; 15'h7E1A: d <= 8'h00; 15'h7E1B: d <= 8'h00;
                15'h7E1C: d <= 8'h00; 15'h7E1D: d <= 8'h00; 15'h7E1E: d <= 8'h00; 15'h7E1F: d <= 8'h00;
                15'h7E20: d <= 8'h00; 15'h7E21: d <= 8'h00; 15'h7E22: d <= 8'h00; 15'h7E23: d <= 8'h00;
                15'h7E24: d <= 8'h00; 15'h7E25: d <= 8'h00; 15'h7E26: d <= 8'h00; 15'h7E27: d <= 8'h00;
                15'h7E28: d <= 8'h00; 15'h7E29: d <= 8'h00; 15'h7E2A: d <= 8'h00; 15'h7E2B: d <= 8'h00;
                15'h7E2C: d <= 8'h00; 15'h7E2D: d <= 8'h00; 15'h7E2E: d <= 8'h00; 15'h7E2F: d <= 8'h7B;
                15'h7E30: d <= 8'h00; 15'h7E31: d <= 8'h00; 15'h7E32: d <= 8'h00; 15'h7E33: d <= 8'h00;
                15'h7E34: d <= 8'h00; 15'h7E35: d <= 8'h00; 15'h7E36: d <= 8'h00; 15'h7E37: d <= 8'h00;
                15'h7E38: d <= 8'h00; 15'h7E39: d <= 8'h00; 15'h7E3A: d <= 8'h00; 15'h7E3B: d <= 8'h00;
                15'h7E3C: d <= 8'h00; 15'h7E3D: d <= 8'h00; 15'h7E3E: d <= 8'h00; 15'h7E3F: d <= 8'h00;
                15'h7E40: d <= 8'h00; 15'h7E41: d <= 8'h00; 15'h7E42: d <= 8'h00; 15'h7E43: d <= 8'h00;
                15'h7E44: d <= 8'h00; 15'h7E45: d <= 8'h00; 15'h7E46: d <= 8'h00; 15'h7E47: d <= 8'h00;
                15'h7E48: d <= 8'h00; 15'h7E49: d <= 8'h00; 15'h7E4A: d <= 8'h00; 15'h7E4B: d <= 8'h00;
                15'h7E4C: d <= 8'h00; 15'h7E4D: d <= 8'h00; 15'h7E4E: d <= 8'h00; 15'h7E4F: d <= 8'h00;
                15'h7E50: d <= 8'h00; 15'h7E51: d <= 8'h00; 15'h7E52: d <= 8'h00; 15'h7E53: d <= 8'h00;
                15'h7E54: d <= 8'h00; 15'h7E55: d <= 8'h00; 15'h7E56: d <= 8'h00; 15'h7E57: d <= 8'h00;
                15'h7E58: d <= 8'h45; 15'h7E59: d <= 8'h35; 15'h7E5A: d <= 8'h32; 15'h7E5B: d <= 8'h00;
                15'h7E5C: d <= 8'h00; 15'h7E5D: d <= 8'h00; 15'h7E5E: d <= 8'h00; 15'h7E5F: d <= 8'h00;
                15'h7E60: d <= 8'h00; 15'h7E61: d <= 8'h00; 15'h7E62: d <= 8'h00; 15'h7E63: d <= 8'h00;
                15'h7E64: d <= 8'h00; 15'h7E65: d <= 8'h00; 15'h7E66: d <= 8'h00; 15'h7E67: d <= 8'h00;
                15'h7E68: d <= 8'h00; 15'h7E69: d <= 8'h00; 15'h7E6A: d <= 8'h00; 15'h7E6B: d <= 8'h00;
                15'h7E6C: d <= 8'h00; 15'h7E6D: d <= 8'h00; 15'h7E6E: d <= 8'h00; 15'h7E6F: d <= 8'h00;
                15'h7E70: d <= 8'h00; 15'h7E71: d <= 8'h00; 15'h7E72: d <= 8'h00; 15'h7E73: d <= 8'h00;
                15'h7E74: d <= 8'h00; 15'h7E75: d <= 8'h00; 15'h7E76: d <= 8'h00; 15'h7E77: d <= 8'h00;
                15'h7E78: d <= 8'h00; 15'h7E79: d <= 8'h00; 15'h7E7A: d <= 8'h00; 15'h7E7B: d <= 8'h00;
                15'h7E7C: d <= 8'h00; 15'h7E7D: d <= 8'h00; 15'h7E7E: d <= 8'h00; 15'h7E7F: d <= 8'hE0;
                15'h7E80: d <= 8'h10; 15'h7E81: d <= 8'h15; 15'h7E82: d <= 8'h1A; 15'h7E83: d <= 8'h1F;
                15'h7E84: d <= 8'h20; 15'h7E85: d <= 8'h25; 15'h7E86: d <= 8'h2A; 15'h7E87: d <= 8'h2F;
                15'h7E88: d <= 8'h34; 15'h7E89: d <= 8'h38; 15'h7E8A: d <= 8'h3C; 15'h7E8B: d <= 8'h31;
                15'h7E8C: d <= 8'h39; 15'h7E8D: d <= 8'h3D; 15'h7E8E: d <= 8'h32; 15'h7E8F: d <= 8'h36;
                15'h7E90: d <= 8'h3E; 15'h7E91: d <= 8'h33; 15'h7E92: d <= 8'h37; 15'h7E93: d <= 8'h3B;
                15'h7E94: d <= 8'h44; 15'h7E95: d <= 8'h48; 15'h7E96: d <= 8'h4C; 15'h7E97: d <= 8'h41;
                15'h7E98: d <= 8'h49; 15'h7E99: d <= 8'h4D; 15'h7E9A: d <= 8'h42; 15'h7E9B: d <= 8'h46;
                15'h7E9C: d <= 8'h4E; 15'h7E9D: d <= 8'h43; 15'h7E9E: d <= 8'h47; 15'h7E9F: d <= 8'h4B;
                15'h7EA0: d <= 8'h50; 15'h7EA1: d <= 8'h55; 15'h7EA2: d <= 8'h5A; 15'h7EA3: d <= 8'h5F;
                15'h7EA4: d <= 8'h60; 15'h7EA5: d <= 8'h65; 15'h7EA6: d <= 8'h6A; 15'h7EA7: d <= 8'h6F;
                15'h7EA8: d <= 8'h74; 15'h7EA9: d <= 8'h78; 15'h7EAA: d <= 8'h7C; 15'h7EAB: d <= 8'h71;
                15'h7EAC: d <= 8'h79; 15'h7EAD: d <= 8'h7D; 15'h7EAE: d <= 8'h72; 15'h7EAF: d <= 8'h76;
                15'h7EB0: d <= 8'h7E; 15'h7EB1: d <= 8'h73; 15'h7EB2: d <= 8'h77; 15'h7EB3: d <= 8'h7B;
                15'h7EB4: d <= 8'h84; 15'h7EB5: d <= 8'h88; 15'h7EB6: d <= 8'h8C; 15'h7EB7: d <= 8'h81;
                15'h7EB8: d <= 8'h89; 15'h7EB9: d <= 8'h8D; 15'h7EBA: d <= 8'h82; 15'h7EBB: d <= 8'h86;
                15'h7EBC: d <= 8'h8E; 15'h7EBD: d <= 8'h83; 15'h7EBE: d <= 8'h87; 15'h7EBF: d <= 8'h8B;
                15'h7EC0: d <= 8'h90; 15'h7EC1: d <= 8'h95; 15'h7EC2: d <= 8'h9A; 15'h7EC3: d <= 8'h9F;
                15'h7EC4: d <= 8'hA4; 15'h7EC5: d <= 8'hA8; 15'h7EC6: d <= 8'hAC; 15'h7EC7: d <= 8'hA1;
                15'h7EC8: d <= 8'hA9; 15'h7EC9: d <= 8'hAD; 15'h7ECA: d <= 8'hA2; 15'h7ECB: d <= 8'hA6;
                15'h7ECC: d <= 8'hAE; 15'h7ECD: d <= 8'hA3; 15'h7ECE: d <= 8'hA7; 15'h7ECF: d <= 8'hAB;
                15'h7ED0: d <= 8'hB4; 15'h7ED1: d <= 8'hB8; 15'h7ED2: d <= 8'hBC; 15'h7ED3: d <= 8'hB1;
                15'h7ED4: d <= 8'hB9; 15'h7ED5: d <= 8'hBD; 15'h7ED6: d <= 8'hB2; 15'h7ED7: d <= 8'hB6;
                15'h7ED8: d <= 8'hBE; 15'h7ED9: d <= 8'hB3; 15'h7EDA: d <= 8'hB7; 15'h7EDB: d <= 8'hBB;
                15'h7EDC: d <= 8'hC4; 15'h7EDD: d <= 8'hC8; 15'h7EDE: d <= 8'hCC; 15'h7EDF: d <= 8'hC1;
                15'h7EE0: d <= 8'hC9; 15'h7EE1: d <= 8'hCD; 15'h7EE2: d <= 8'hC2; 15'h7EE3: d <= 8'hC6;
                15'h7EE4: d <= 8'hCE; 15'h7EE5: d <= 8'hC3; 15'h7EE6: d <= 8'hC7; 15'h7EE7: d <= 8'hCB;
                15'h7EE8: d <= 8'hC0; 15'h7EE9: d <= 8'hC5; 15'h7EEA: d <= 8'hCA; 15'h7EEB: d <= 8'hCF;
                15'h7EEC: d <= 8'hD0; 15'h7EED: d <= 8'hD5; 15'h7EEE: d <= 8'hDA; 15'h7EEF: d <= 8'hDF;
                15'h7EF0: d <= 8'h74; 15'h7EF1: d <= 8'h78; 15'h7EF2: d <= 8'h7C; 15'h7EF3: d <= 8'h71;
                15'h7EF4: d <= 8'h79; 15'h7EF5: d <= 8'h7D; 15'h7EF6: d <= 8'h72; 15'h7EF7: d <= 8'h76;
                15'h7EF8: d <= 8'h7E; 15'h7EF9: d <= 8'h73; 15'h7EFA: d <= 8'h77; 15'h7EFB: d <= 8'h7B;
                15'h7EFC: d <= 8'hA0; 15'h7EFD: d <= 8'hA5; 15'h7EFE: d <= 8'hAA; 15'h7EFF: d <= 8'hAF;
                15'h7F00: d <= 8'h00; 15'h7F01: d <= 8'h00; 15'h7F02: d <= 8'h00; 15'h7F03: d <= 8'h00;
                15'h7F04: d <= 8'h00; 15'h7F05: d <= 8'h00; 15'h7F06: d <= 8'h00; 15'h7F07: d <= 8'h00;
                15'h7F08: d <= 8'h00; 15'h7F09: d <= 8'h00; 15'h7F0A: d <= 8'h00; 15'h7F0B: d <= 8'h00;
                15'h7F0C: d <= 8'h00; 15'h7F0D: d <= 8'h00; 15'h7F0E: d <= 8'h00; 15'h7F0F: d <= 8'h00;
                15'h7F10: d <= 8'h00; 15'h7F11: d <= 8'h00; 15'h7F12: d <= 8'h00; 15'h7F13: d <= 8'h00;
                15'h7F14: d <= 8'h00; 15'h7F15: d <= 8'h00; 15'h7F16: d <= 8'h00; 15'h7F17: d <= 8'h00;
                15'h7F18: d <= 8'h00; 15'h7F19: d <= 8'h00; 15'h7F1A: d <= 8'h00; 15'h7F1B: d <= 8'h00;
                15'h7F1C: d <= 8'h00; 15'h7F1D: d <= 8'h00; 15'h7F1E: d <= 8'h00; 15'h7F1F: d <= 8'h00;
                15'h7F20: d <= 8'h00; 15'h7F21: d <= 8'h00; 15'h7F22: d <= 8'h00; 15'h7F23: d <= 8'h00;
                15'h7F24: d <= 8'h00; 15'h7F25: d <= 8'h00; 15'h7F26: d <= 8'h00; 15'h7F27: d <= 8'h00;
                15'h7F28: d <= 8'h00; 15'h7F29: d <= 8'h00; 15'h7F2A: d <= 8'h00; 15'h7F2B: d <= 8'h00;
                15'h7F2C: d <= 8'h00; 15'h7F2D: d <= 8'h00; 15'h7F2E: d <= 8'h00; 15'h7F2F: d <= 8'h7B;
                15'h7F30: d <= 8'h00; 15'h7F31: d <= 8'h00; 15'h7F32: d <= 8'h00; 15'h7F33: d <= 8'h00;
                15'h7F34: d <= 8'h00; 15'h7F35: d <= 8'h00; 15'h7F36: d <= 8'h00; 15'h7F37: d <= 8'h00;
                15'h7F38: d <= 8'h00; 15'h7F39: d <= 8'h00; 15'h7F3A: d <= 8'h00; 15'h7F3B: d <= 8'h00;
                15'h7F3C: d <= 8'h00; 15'h7F3D: d <= 8'h00; 15'h7F3E: d <= 8'h00; 15'h7F3F: d <= 8'h00;
                15'h7F40: d <= 8'h00; 15'h7F41: d <= 8'h00; 15'h7F42: d <= 8'h00; 15'h7F43: d <= 8'h00;
                15'h7F44: d <= 8'h00; 15'h7F45: d <= 8'h00; 15'h7F46: d <= 8'h00; 15'h7F47: d <= 8'h00;
                15'h7F48: d <= 8'h00; 15'h7F49: d <= 8'h00; 15'h7F4A: d <= 8'h00; 15'h7F4B: d <= 8'h00;
                15'h7F4C: d <= 8'h00; 15'h7F4D: d <= 8'h00; 15'h7F4E: d <= 8'h00; 15'h7F4F: d <= 8'h00;
                15'h7F50: d <= 8'h00; 15'h7F51: d <= 8'h00; 15'h7F52: d <= 8'h00; 15'h7F53: d <= 8'h00;
                15'h7F54: d <= 8'h00; 15'h7F55: d <= 8'h00; 15'h7F56: d <= 8'h00; 15'h7F57: d <= 8'h00;
                15'h7F58: d <= 8'h45; 15'h7F59: d <= 8'h35; 15'h7F5A: d <= 8'h32; 15'h7F5B: d <= 8'h00;
                15'h7F5C: d <= 8'h00; 15'h7F5D: d <= 8'h00; 15'h7F5E: d <= 8'h00; 15'h7F5F: d <= 8'h00;
                15'h7F60: d <= 8'h00; 15'h7F61: d <= 8'h00; 15'h7F62: d <= 8'h00; 15'h7F63: d <= 8'h00;
                15'h7F64: d <= 8'h00; 15'h7F65: d <= 8'h00; 15'h7F66: d <= 8'h00; 15'h7F67: d <= 8'h00;
                15'h7F68: d <= 8'h00; 15'h7F69: d <= 8'h00; 15'h7F6A: d <= 8'h00; 15'h7F6B: d <= 8'h00;
                15'h7F6C: d <= 8'h00; 15'h7F6D: d <= 8'h00; 15'h7F6E: d <= 8'h00; 15'h7F6F: d <= 8'h00;
                15'h7F70: d <= 8'h00; 15'h7F71: d <= 8'h00; 15'h7F72: d <= 8'h00; 15'h7F73: d <= 8'h00;
                15'h7F74: d <= 8'h00; 15'h7F75: d <= 8'h00; 15'h7F76: d <= 8'h00; 15'h7F77: d <= 8'h00;
                15'h7F78: d <= 8'h00; 15'h7F79: d <= 8'h00; 15'h7F7A: d <= 8'h00; 15'h7F7B: d <= 8'h00;
                15'h7F7C: d <= 8'h00; 15'h7F7D: d <= 8'h00; 15'h7F7E: d <= 8'h00; 15'h7F7F: d <= 8'hE0;
                15'h7F80: d <= 8'h10; 15'h7F81: d <= 8'h15; 15'h7F82: d <= 8'h1A; 15'h7F83: d <= 8'h1F;
                15'h7F84: d <= 8'h20; 15'h7F85: d <= 8'h25; 15'h7F86: d <= 8'h2A; 15'h7F87: d <= 8'h2F;
                15'h7F88: d <= 8'h34; 15'h7F89: d <= 8'h38; 15'h7F8A: d <= 8'h3C; 15'h7F8B: d <= 8'h31;
                15'h7F8C: d <= 8'h39; 15'h7F8D: d <= 8'h3D; 15'h7F8E: d <= 8'h32; 15'h7F8F: d <= 8'h36;
                15'h7F90: d <= 8'h3E; 15'h7F91: d <= 8'h33; 15'h7F92: d <= 8'h37; 15'h7F93: d <= 8'h3B;
                15'h7F94: d <= 8'h44; 15'h7F95: d <= 8'h48; 15'h7F96: d <= 8'h4C; 15'h7F97: d <= 8'h41;
                15'h7F98: d <= 8'h49; 15'h7F99: d <= 8'h4D; 15'h7F9A: d <= 8'h42; 15'h7F9B: d <= 8'h46;
                15'h7F9C: d <= 8'h4E; 15'h7F9D: d <= 8'h43; 15'h7F9E: d <= 8'h47; 15'h7F9F: d <= 8'h4B;
                15'h7FA0: d <= 8'h50; 15'h7FA1: d <= 8'h55; 15'h7FA2: d <= 8'h5A; 15'h7FA3: d <= 8'h5F;
                15'h7FA4: d <= 8'h60; 15'h7FA5: d <= 8'h65; 15'h7FA6: d <= 8'h6A; 15'h7FA7: d <= 8'h6F;
                15'h7FA8: d <= 8'h74; 15'h7FA9: d <= 8'h78; 15'h7FAA: d <= 8'h7C; 15'h7FAB: d <= 8'h71;
                15'h7FAC: d <= 8'h79; 15'h7FAD: d <= 8'h7D; 15'h7FAE: d <= 8'h72; 15'h7FAF: d <= 8'h76;
                15'h7FB0: d <= 8'h7E; 15'h7FB1: d <= 8'h73; 15'h7FB2: d <= 8'h77; 15'h7FB3: d <= 8'h7B;
                15'h7FB4: d <= 8'h84; 15'h7FB5: d <= 8'h88; 15'h7FB6: d <= 8'h8C; 15'h7FB7: d <= 8'h81;
                15'h7FB8: d <= 8'h89; 15'h7FB9: d <= 8'h8D; 15'h7FBA: d <= 8'h82; 15'h7FBB: d <= 8'h86;
                15'h7FBC: d <= 8'h8E; 15'h7FBD: d <= 8'h83; 15'h7FBE: d <= 8'h87; 15'h7FBF: d <= 8'h8B;
                15'h7FC0: d <= 8'h90; 15'h7FC1: d <= 8'h95; 15'h7FC2: d <= 8'h9A; 15'h7FC3: d <= 8'h9F;
                15'h7FC4: d <= 8'hA4; 15'h7FC5: d <= 8'hA8; 15'h7FC6: d <= 8'hAC; 15'h7FC7: d <= 8'hA1;
                15'h7FC8: d <= 8'hA9; 15'h7FC9: d <= 8'hAD; 15'h7FCA: d <= 8'hA2; 15'h7FCB: d <= 8'hA6;
                15'h7FCC: d <= 8'hAE; 15'h7FCD: d <= 8'hA3; 15'h7FCE: d <= 8'hA7; 15'h7FCF: d <= 8'hAB;
                15'h7FD0: d <= 8'hB4; 15'h7FD1: d <= 8'hB8; 15'h7FD2: d <= 8'hBC; 15'h7FD3: d <= 8'hB1;
                15'h7FD4: d <= 8'hB9; 15'h7FD5: d <= 8'hBD; 15'h7FD6: d <= 8'hB2; 15'h7FD7: d <= 8'hB6;
                15'h7FD8: d <= 8'hBE; 15'h7FD9: d <= 8'hB3; 15'h7FDA: d <= 8'hB7; 15'h7FDB: d <= 8'hBB;
                15'h7FDC: d <= 8'hC4; 15'h7FDD: d <= 8'hC8; 15'h7FDE: d <= 8'hCC; 15'h7FDF: d <= 8'hC1;
                15'h7FE0: d <= 8'hC9; 15'h7FE1: d <= 8'hCD; 15'h7FE2: d <= 8'hC2; 15'h7FE3: d <= 8'hC6;
                15'h7FE4: d <= 8'hCE; 15'h7FE5: d <= 8'hC3; 15'h7FE6: d <= 8'hC7; 15'h7FE7: d <= 8'hCB;
                15'h7FE8: d <= 8'hC0; 15'h7FE9: d <= 8'hC5; 15'h7FEA: d <= 8'hCA; 15'h7FEB: d <= 8'hCF;
                15'h7FEC: d <= 8'hD0; 15'h7FED: d <= 8'hD5; 15'h7FEE: d <= 8'hDA; 15'h7FEF: d <= 8'hDF;
                15'h7FF0: d <= 8'h74; 15'h7FF1: d <= 8'h78; 15'h7FF2: d <= 8'h7C; 15'h7FF3: d <= 8'h71;
                15'h7FF4: d <= 8'h79; 15'h7FF5: d <= 8'h7D; 15'h7FF6: d <= 8'h72; 15'h7FF7: d <= 8'h76;
                15'h7FF8: d <= 8'h7E; 15'h7FF9: d <= 8'h73; 15'h7FFA: d <= 8'h77; 15'h7FFB: d <= 8'h7B;
                15'h7FFC: d <= 8'hA0; 15'h7FFD: d <= 8'hA5; 15'h7FFE: d <= 8'hAA; 15'h7FFF: d <= 8'hAF;
                            endcase
    end //end:always_posedge_clk
    assign dout = d;
endmodule //end:pipeline_rom_1a
