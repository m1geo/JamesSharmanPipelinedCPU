// -----------------------------------------------------------------------------
// Title   : Memory (RAM & ROM) (MainBus/memory.v)
// Create  : Tue 20 Dec 22:32:02 GMT 2022
//
// Name    : JAM-1 8-bit Pipelined CPU in Verilog
// Author  : George Smart, M1GEO.  https://www.george-smart.co.uk
// GitHub  : https://github.com/m1geo/JamesSharmanPipelinedCPU
// CPU Dsn : James Sharman; Video Series => https://youtu.be/3iHag4k4yEg
//
// Desc.   : Combined RAM+ROM to use BRAM in FPGA
// -----------------------------------------------------------------------------

module memory
(
    // ports here
);

    // code here

endmodule //end:memory
