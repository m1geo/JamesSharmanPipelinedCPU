/*

Name:				ALU?
Schematic Source:   ??
Schematic Rev:		??
Designer:			James Sharman (weirdboyjim)

FPGA/Verilog: 		George Smart (@m1geo) http://www.george-smart.co.uk
Project Source:		https://github.com/m1geo/JamesSharmanPipelinedCPU

Module notes:
	See video part 34, diagram at 32 seconds: https://www.youtube.com/watch?v=pMV_0qT0uY0?t=32
	The entire ALU is shown.
	Verilog is missing for "ADD", "FLAGS" and "ZERO CMP".
*/

module ALU ();

	// main code goes here!

endmodule